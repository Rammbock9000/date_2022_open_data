--------------------------------------------------------------------------------
--                         ModuloCounter_14_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_14_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of ModuloCounter_14_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(3 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 13 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_5_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_5_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(2 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_5_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000",
         iS_1 when "001",
         iS_2 when "010",
         iS_3 when "011",
         iS_4 when "100",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid2513963_RightShifter
--                (RightShifter_24_by_max_26_F250_uid2513965)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2513963_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2513963_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid2513968
--                  (IntAdderAlternative_27_f250_uid2513972)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid2513968 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid2513968 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid2513975
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid2513975 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid2513975 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid2513978
--                   (IntAdderClassical_34_f250_uid2513980)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid2513978 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid2513978 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid2513963
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2513963 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2513963 is
   component FPAdd_8_23_uid2513963_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid2513968 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid2513975 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid2513978 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid2513963_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid2513968  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid2513975  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid2513978  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid2513963 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid2513963  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_14_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_14_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_14_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
         iS_9 when "1001",
         iS_10 when "1010",
         iS_11 when "1011",
         iS_12 when "1100",
         iS_13 when "1101",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2515284
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2515284 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2515284 is
signal XX_m2515285 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m2515285 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m2515285 <= X ;
   YY_m2515285 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_33_f500_uid2515288
--                   (IntAdderClassical_33_f500_uid2515290)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid2515288 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid2515288 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2515284 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid2515288 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2515284  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
      RoundingAdder: IntAdder_33_f500_uid2515288  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid2515547_RightShifter
--                (RightShifter_24_by_max_26_F250_uid2515549)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2515547_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2515547_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid2515552
--                  (IntAdderAlternative_27_f250_uid2515556)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid2515552 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid2515552 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid2515559
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid2515559 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid2515559 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid2515562
--                   (IntAdderClassical_34_f250_uid2515564)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid2515562 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid2515562 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid2515547
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2515547 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2515547 is
   component FPAdd_8_23_uid2515547_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid2515552 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid2515559 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid2515562 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid2515547_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid2515552  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid2515559  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid2515562  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   component FPAdd_8_23_uid2515547 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= (Y(Y'length-1 downto Y'length-2)) & (not Y(Y'length-3)) & Y(Y'length-4 downto 0);
   FPAddSubOp_instance: FPAdd_8_23_uid2515547  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_13_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_13_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_13_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
         iS_9 when "1001",
         iS_10 when "1010",
         iS_11 when "1011",
         iS_12 when "1100",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_9_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_9_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_9_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_0_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_0_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_0_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_2_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_2_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_2_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn5_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn5_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn5_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn3_mult_pi_div_4_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn3_mult_pi_div_4_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn3_mult_pi_div_4_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111001101010000010011110011";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_cosn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--             Constant_float_8_23_sinn7_mult_pi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinn7_mult_pi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinn7_mult_pi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_cosnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_cosnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_cosnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111011011001000001101011110";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_sinnpi_div_8_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_sinnpi_div_8_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_sinnpi_div_8_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111110110000111110111100010101";
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      Y <= s11;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      Y <= s10;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      Y <= s9;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      Y <= s7;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      Y <= s12;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "000" when "0001",
      "000" when "0010",
      "001" when "0011",
      "000" when "0100",
      "000" when "0101",
      "010" when "0110",
      "000" when "0111",
      "000" when "1000",
      "011" when "1001",
      "000" when "1010",
      "100" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "001" when "0100",
      "000" when "0101",
      "000" when "0110",
      "010" when "0111",
      "000" when "1000",
      "000" when "1001",
      "011" when "1010",
      "000" when "1011",
      "100" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "001" when "0110",
      "000" when "0111",
      "000" when "1000",
      "010" when "1001",
      "000" when "1010",
      "000" when "1011",
      "011" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "100" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "000" when "1001",
      "010" when "1010",
      "000" when "1011",
      "000" when "1100",
      "011" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "001" when "0001",
      "000" when "0010",
      "000" when "0011",
      "010" when "0100",
      "000" when "0101",
      "000" when "0110",
      "011" when "0111",
      "000" when "1000",
      "100" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "001" when "0001",
      "000" when "0010",
      "000" when "0011",
      "010" when "0100",
      "000" when "0101",
      "000" when "0110",
      "011" when "0111",
      "000" when "1000",
      "100" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "011" when "0000",
      "000" when "0001",
      "100" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "000" when "0111",
      "001" when "1000",
      "000" when "1001",
      "000" when "1010",
      "010" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "011" when "0000",
      "000" when "0001",
      "100" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "000" when "0111",
      "001" when "1000",
      "000" when "1001",
      "000" when "1010",
      "010" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "001" when "0100",
      "000" when "0101",
      "000" when "0110",
      "010" when "0111",
      "000" when "1000",
      "000" when "1001",
      "011" when "1010",
      "000" when "1011",
      "100" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "001" when "0100",
      "000" when "0101",
      "000" when "0110",
      "010" when "0111",
      "000" when "1000",
      "000" when "1001",
      "011" when "1010",
      "000" when "1011",
      "100" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "100" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "000" when "1001",
      "010" when "1010",
      "000" when "1011",
      "000" when "1100",
      "011" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "100" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "000" when "1001",
      "010" when "1010",
      "000" when "1011",
      "000" when "1100",
      "011" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "000" when "0001",
      "000" when "0010",
      "001" when "0011",
      "000" when "0100",
      "000" when "0101",
      "010" when "0110",
      "000" when "0111",
      "000" when "1000",
      "011" when "1001",
      "000" when "1010",
      "100" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "000" when "0001",
      "000" when "0010",
      "001" when "0011",
      "000" when "0100",
      "000" when "0101",
      "010" when "0110",
      "000" when "0111",
      "000" when "1000",
      "011" when "1001",
      "000" when "1010",
      "100" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "100" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "000" when "1001",
      "010" when "1010",
      "000" when "1011",
      "000" when "1100",
      "011" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "011" when "0000",
      "000" when "0001",
      "100" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "000" when "0111",
      "001" when "1000",
      "000" when "1001",
      "000" when "1010",
      "010" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "000" when "0001",
      "000" when "0010",
      "001" when "0011",
      "000" when "0100",
      "000" when "0101",
      "010" when "0110",
      "000" when "0111",
      "000" when "1000",
      "011" when "1001",
      "000" when "1010",
      "100" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "000" when "0001",
      "000" when "0010",
      "001" when "0011",
      "000" when "0100",
      "000" when "0101",
      "010" when "0110",
      "000" when "0111",
      "000" when "1000",
      "011" when "1001",
      "000" when "1010",
      "100" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "001" when "0110",
      "000" when "0111",
      "000" when "1000",
      "010" when "1001",
      "000" when "1010",
      "000" when "1011",
      "011" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "100" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "001" when "0110",
      "000" when "0111",
      "000" when "1000",
      "010" when "1001",
      "000" when "1010",
      "000" when "1011",
      "011" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "001" when "0001",
      "000" when "0010",
      "000" when "0011",
      "010" when "0100",
      "000" when "0101",
      "000" when "0110",
      "011" when "0111",
      "000" when "1000",
      "100" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "001" when "0001",
      "000" when "0010",
      "000" when "0011",
      "010" when "0100",
      "000" when "0101",
      "000" when "0110",
      "011" when "0111",
      "000" when "1000",
      "100" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "011" when "0000",
      "000" when "0001",
      "100" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "000" when "0111",
      "001" when "1000",
      "000" when "1001",
      "000" when "1010",
      "010" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "011" when "0000",
      "000" when "0001",
      "100" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "000" when "0111",
      "001" when "1000",
      "000" when "1001",
      "000" when "1010",
      "010" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "001" when "0100",
      "000" when "0101",
      "000" when "0110",
      "010" when "0111",
      "000" when "1000",
      "000" when "1001",
      "011" when "1010",
      "000" when "1011",
      "100" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "000" when "0001",
      "000" when "0010",
      "000" when "0011",
      "001" when "0100",
      "000" when "0101",
      "000" when "0110",
      "010" when "0111",
      "000" when "1000",
      "000" when "1001",
      "011" when "1010",
      "000" when "1011",
      "100" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "100" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "000" when "1001",
      "010" when "1010",
      "000" when "1011",
      "000" when "1100",
      "011" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "100" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "000" when "1001",
      "010" when "1010",
      "000" when "1011",
      "000" when "1100",
      "011" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "001" when "0001",
      "000" when "0010",
      "000" when "0011",
      "010" when "0100",
      "000" when "0101",
      "000" when "0110",
      "011" when "0111",
      "000" when "1000",
      "100" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "001" when "0001",
      "000" when "0010",
      "000" when "0011",
      "010" when "0100",
      "000" when "0101",
      "000" when "0110",
      "011" when "0111",
      "000" when "1000",
      "100" when "1001",
      "000" when "1010",
      "000" when "1011",
      "000" when "1100",
      "000" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "100" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "000" when "1001",
      "010" when "1010",
      "000" when "1011",
      "000" when "1100",
      "011" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--             GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "100" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "000" when "0101",
      "000" when "0110",
      "001" when "0111",
      "000" when "1000",
      "000" when "1001",
      "010" when "1010",
      "000" when "1011",
      "000" when "1100",
      "011" when "1101",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--    GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product326_4_impl_0_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product326_4_impl_0_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product326_4_impl_0_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0011" when "0000",
      "0111" when "0001",
      "0010" when "0010",
      "1011" when "0011",
      "1100" when "0100",
      "0000" when "0101",
      "1010" when "0110",
      "1000" when "0111",
      "0000" when "1000",
      "0001" when "1001",
      "0110" when "1010",
      "1001" when "1011",
      "0101" when "1100",
      "0100" when "1101",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product326_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product326_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product326_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product326_4_impl_0_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product326_4_impl_0_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product326_4_impl_1_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product326_4_impl_1_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product326_4_impl_1_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "1011" when "0000",
      "0110" when "0001",
      "1010" when "0010",
      "0011" when "0011",
      "0100" when "0100",
      "1100" when "0101",
      "0010" when "0110",
      "0000" when "0111",
      "0000" when "1000",
      "1001" when "1001",
      "1000" when "1010",
      "0001" when "1011",
      "0111" when "1100",
      "0101" when "1101",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product326_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product326_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product326_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product326_4_impl_1_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product326_4_impl_1_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product237_4_impl_0_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product237_4_impl_0_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product237_4_impl_0_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0000" when "0000",
      "0100" when "0001",
      "0000" when "0010",
      "1000" when "0011",
      "0000" when "0100",
      "0000" when "0101",
      "0111" when "0110",
      "0101" when "0111",
      "0000" when "1000",
      "0110" when "1001",
      "0010" when "1010",
      "0000" when "1011",
      "0001" when "1100",
      "0011" when "1101",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product237_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product237_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product237_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product237_4_impl_0_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product237_4_impl_0_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product237_4_impl_1_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product237_4_impl_1_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product237_4_impl_1_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0000" when "0000",
      "0100" when "0001",
      "0000" when "0010",
      "0011" when "0011",
      "1000" when "0100",
      "0000" when "0101",
      "0010" when "0110",
      "0000" when "0111",
      "0000" when "1000",
      "0001" when "1001",
      "0111" when "1010",
      "0000" when "1011",
      "0110" when "1100",
      "0101" when "1101",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product237_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product237_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product237_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product237_4_impl_1_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product237_4_impl_1_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 23 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      Y <= s22;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 15 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      Y <= s14;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      Y <= s13;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 17 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      Y <= s16;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 16 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      Y <= s15;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      Y <= s20;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 20 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      Y <= s19;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      Y <= s8;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 22 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      Y <= s21;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          x0_re_0 : in std_logic_vector(31 downto 0);
          x0_im_0 : in std_logic_vector(31 downto 0);
          x1_re_0 : in std_logic_vector(31 downto 0);
          x1_im_0 : in std_logic_vector(31 downto 0);
          x2_re_0 : in std_logic_vector(31 downto 0);
          x2_im_0 : in std_logic_vector(31 downto 0);
          x3_re_0 : in std_logic_vector(31 downto 0);
          x3_im_0 : in std_logic_vector(31 downto 0);
          x4_re_0 : in std_logic_vector(31 downto 0);
          x4_im_0 : in std_logic_vector(31 downto 0);
          x5_re_0 : in std_logic_vector(31 downto 0);
          x5_im_0 : in std_logic_vector(31 downto 0);
          x6_re_0 : in std_logic_vector(31 downto 0);
          x6_im_0 : in std_logic_vector(31 downto 0);
          x7_re_0 : in std_logic_vector(31 downto 0);
          x7_im_0 : in std_logic_vector(31 downto 0);
          x8_re_0 : in std_logic_vector(31 downto 0);
          x8_im_0 : in std_logic_vector(31 downto 0);
          x9_re_0 : in std_logic_vector(31 downto 0);
          x9_im_0 : in std_logic_vector(31 downto 0);
          x10_re_0 : in std_logic_vector(31 downto 0);
          x10_im_0 : in std_logic_vector(31 downto 0);
          x11_re_0 : in std_logic_vector(31 downto 0);
          x11_im_0 : in std_logic_vector(31 downto 0);
          x12_re_0 : in std_logic_vector(31 downto 0);
          x12_im_0 : in std_logic_vector(31 downto 0);
          x13_re_0 : in std_logic_vector(31 downto 0);
          x13_im_0 : in std_logic_vector(31 downto 0);
          x14_re_0 : in std_logic_vector(31 downto 0);
          x14_im_0 : in std_logic_vector(31 downto 0);
          x15_re_0 : in std_logic_vector(31 downto 0);
          x15_im_0 : in std_logic_vector(31 downto 0);
          y0_re_0 : out std_logic_vector(31 downto 0);
          y0_im_0 : out std_logic_vector(31 downto 0);
          y1_re_0 : out std_logic_vector(31 downto 0);
          y1_im_0 : out std_logic_vector(31 downto 0);
          y2_re_0 : out std_logic_vector(31 downto 0);
          y2_im_0 : out std_logic_vector(31 downto 0);
          y3_re_0 : out std_logic_vector(31 downto 0);
          y3_im_0 : out std_logic_vector(31 downto 0);
          y4_re_0 : out std_logic_vector(31 downto 0);
          y4_im_0 : out std_logic_vector(31 downto 0);
          y5_re_0 : out std_logic_vector(31 downto 0);
          y5_im_0 : out std_logic_vector(31 downto 0);
          y6_re_0 : out std_logic_vector(31 downto 0);
          y6_im_0 : out std_logic_vector(31 downto 0);
          y7_re_0 : out std_logic_vector(31 downto 0);
          y7_im_0 : out std_logic_vector(31 downto 0);
          y8_re_0 : out std_logic_vector(31 downto 0);
          y8_im_0 : out std_logic_vector(31 downto 0);
          y9_re_0 : out std_logic_vector(31 downto 0);
          y9_im_0 : out std_logic_vector(31 downto 0);
          y10_re_0 : out std_logic_vector(31 downto 0);
          y10_im_0 : out std_logic_vector(31 downto 0);
          y11_re_0 : out std_logic_vector(31 downto 0);
          y11_im_0 : out std_logic_vector(31 downto 0);
          y12_re_0 : out std_logic_vector(31 downto 0);
          y12_im_0 : out std_logic_vector(31 downto 0);
          y13_re_0 : out std_logic_vector(31 downto 0);
          y13_im_0 : out std_logic_vector(31 downto 0);
          y14_re_0 : out std_logic_vector(31 downto 0);
          y14_im_0 : out std_logic_vector(31 downto 0);
          y15_re_0 : out std_logic_vector(31 downto 0);
          y15_im_0 : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_14_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(3 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_5_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(2 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_14_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_13_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_9_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_0_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_2_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn5_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn3_mult_pi_div_4_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinn7_mult_pi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_cosnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_sinnpi_div_8_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product326_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product326_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product237_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product237_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount141_out : std_logic_vector(3 downto 0) := (others => '0');
signal x0_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x1_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x2_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x3_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x4_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x5_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x6_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x7_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x8_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x9_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x10_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x11_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x12_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x13_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x14_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_re_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal x15_im_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y1_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y1_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y2_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y2_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y3_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y3_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y4_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y4_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y5_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y5_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y6_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y6_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y7_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y7_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y8_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y8_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y9_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y9_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y10_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y10_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y11_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y11_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y12_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y12_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y13_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y13_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y14_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y14_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y15_re_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y15_im_0_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add2_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add2_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add11_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add11_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add3_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add3_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add12_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add12_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add9_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add9_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add9_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add9_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add9_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add18_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add18_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add18_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add18_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add18_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add18_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add128_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add128_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add128_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add128_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add128_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add128_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add40_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add40_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add40_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add40_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add40_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add40_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product4_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product4_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product11_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product11_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product21_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product21_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product31_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product31_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract2_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract2_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product5_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product5_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product5_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product5_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product5_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product5_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product12_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product12_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product22_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product22_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product32_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product32_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product6_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product6_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No200_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No201_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No202_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No203_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product23_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No204_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product23_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No205_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No206_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No207_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No208_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No209_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No210_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No211_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No212_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No213_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product33_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No214_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product33_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract4_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract4_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product37_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product37_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product37_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product37_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product37_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product37_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract9_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract9_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product39_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product39_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product39_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract20_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract20_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract20_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract20_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No254_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No255_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract20_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No256_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract20_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No257_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product220_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product220_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No258_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product220_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No259_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product220_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product220_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No260_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product220_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No261_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product220_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product220_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No262_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product220_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No263_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product323_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No264_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No265_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product323_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No266_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No267_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product323_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No268_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No269_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product323_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No270_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product323_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No271_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product325_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product325_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No272_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product325_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No273_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product325_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product325_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No274_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product325_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No275_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract26_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No276_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No277_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract26_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No278_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No279_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract26_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No280_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No281_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract26_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No282_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No283_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract26_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No284_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract26_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No285_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product55_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No286_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No287_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product55_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No288_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No289_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product55_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No290_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product55_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No291_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product226_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No292_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No293_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product226_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No294_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product226_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No295_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product326_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product326_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No296_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product326_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No297_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract29_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract29_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No298_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract29_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No299_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract29_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract29_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No300_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract29_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No301_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract29_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract29_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No302_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract29_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No303_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract29_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract29_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No304_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract29_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No305_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract29_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract29_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No306_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract29_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No307_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract33_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract33_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No308_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract33_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No309_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract33_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract33_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No310_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract33_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No311_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract33_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract33_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No312_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract33_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No313_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract33_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract33_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No314_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract33_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No315_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract33_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract33_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No316_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract33_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No317_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product237_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product237_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No318_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product237_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No319_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract38_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract38_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No320_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract38_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No321_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract38_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract38_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No322_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract38_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No323_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract38_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract38_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No324_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract38_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No325_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract38_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract38_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No326_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract38_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No327_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract38_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract38_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No328_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract38_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No329_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant13_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant5_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant14_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant15_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant7_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant16_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant8_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant17_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant18_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No206_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No214_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay28No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay28No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay28No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay28No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay28No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No249_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No252_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_y0_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y0_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y1_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y1_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y2_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y2_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y3_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y3_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y4_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y4_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y5_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y5_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y6_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y6_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y7_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y7_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y8_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y8_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y9_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y9_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y10_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y10_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y11_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y11_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y12_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y12_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y13_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y13_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y14_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y14_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y15_re_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_y15_im_0_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Product326_4_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product326_4_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product237_4_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product237_4_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out : std_logic_vector(33 downto 0) := (others => '0');
signal x0_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x0_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x1_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x2_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x3_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x4_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x5_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x6_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x7_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x8_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x9_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x10_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x11_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x12_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x13_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x14_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal x15_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal y0_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y0_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y1_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y1_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y2_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y2_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y3_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y3_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y4_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y4_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y5_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y5_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y6_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y6_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y7_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y7_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y8_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y8_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y9_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y9_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y10_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y10_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y11_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y11_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y12_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y12_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y13_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y13_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y14_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y14_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y15_re_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal y15_im_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out_to_Add3_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out_to_Add3_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out_to_Add3_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out_to_Add3_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out_to_Add3_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out_to_Add3_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out_to_Add3_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out_to_Add3_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out_to_Add3_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out_to_Add3_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out_to_Add12_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out_to_Add12_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No60_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No75_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No20_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay28No_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out_to_Add12_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out_to_Add12_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No61_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No76_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No21_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay28No1_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out_to_Add12_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out_to_Add12_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No62_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No22_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay28No2_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out_to_Add12_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out_to_Add12_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No63_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No23_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay28No3_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out_to_Add12_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out_to_Add12_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No64_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No24_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay28No4_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out_to_Add9_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out_to_Add9_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No15_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out_to_Add9_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out_to_Add9_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No16_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out_to_Add9_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out_to_Add9_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No17_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out_to_Add9_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out_to_Add9_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No18_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out_to_Add9_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out_to_Add9_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay27No19_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out_to_Add18_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out_to_Add18_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No10_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out_to_Add18_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out_to_Add18_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No11_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out_to_Add18_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out_to_Add18_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No12_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out_to_Add18_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out_to_Add18_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No13_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out_to_Add18_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out_to_Add18_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No14_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out_to_Add128_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out_to_Add128_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No25_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out_to_Add128_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out_to_Add128_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No71_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No26_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out_to_Add128_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out_to_Add128_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No27_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out_to_Add128_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out_to_Add128_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No28_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out_to_Add128_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out_to_Add128_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay4No74_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No214_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No29_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out_to_Add40_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out_to_Add40_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No30_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No35_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out_to_Add40_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out_to_Add40_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No31_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No1_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No36_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out_to_Add40_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out_to_Add40_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No2_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No32_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No37_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No252_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out_to_Add40_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out_to_Add40_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No33_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No3_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No38_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out_to_Add40_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out_to_Add40_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay11No34_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No4_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No39_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No1_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No2_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out_to_Product11_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out_to_Product11_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out_to_Product11_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out_to_Product11_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No4_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No4_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out_to_Product21_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out_to_Product21_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out_to_Product21_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out_to_Product21_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No3_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out_to_Product31_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out_to_Product31_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No1_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out_to_Product31_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out_to_Product31_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No10_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No25_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No11_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No26_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No12_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No42_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No27_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No43_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No28_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No13_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No14_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No29_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out_to_Product5_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out_to_Product5_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out_to_Product5_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out_to_Product5_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out_to_Product5_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out_to_Product5_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay10No2_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out_to_Product5_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out_to_Product5_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out_to_Product5_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out_to_Product5_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out_to_Product12_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out_to_Product12_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out_to_Product12_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out_to_Product12_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out_to_Product12_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out_to_Product12_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out_to_Product12_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out_to_Product12_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out_to_Product12_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out_to_Product12_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out_to_Product22_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out_to_Product22_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out_to_Product22_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out_to_Product22_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out_to_Product22_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out_to_Product22_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out_to_Product22_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out_to_Product22_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out_to_Product22_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out_to_Product22_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out_to_Product32_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out_to_Product32_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out_to_Product6_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out_to_Product6_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out_to_Product6_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out_to_Product6_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out_to_Product6_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out_to_Product6_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out_to_Product6_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out_to_Product6_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out_to_Product6_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out_to_Product6_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out_to_Product23_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out_to_Product23_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out_to_Product23_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out_to_Product23_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No200_out_to_Product23_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No201_out_to_Product23_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No202_out_to_Product23_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No203_out_to_Product23_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No204_out_to_Product23_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No205_out_to_Product23_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No206_out_to_Product33_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No207_out_to_Product33_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No208_out_to_Product33_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No209_out_to_Product33_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No210_out_to_Product33_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No211_out_to_Product33_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No212_out_to_Product33_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No213_out_to_Product33_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No214_out_to_Product33_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out_to_Product33_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out_to_Subtract4_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out_to_Subtract4_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No15_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No5_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out_to_Subtract4_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out_to_Subtract4_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No16_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No6_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out_to_Subtract4_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out_to_Subtract4_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No17_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No7_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out_to_Subtract4_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out_to_Subtract4_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No18_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No8_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out_to_Subtract4_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out_to_Subtract4_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No19_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay16No9_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out_to_Product37_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out_to_Product37_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out_to_Product37_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out_to_Product37_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out_to_Product37_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out_to_Product37_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out_to_Product37_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out_to_Product37_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out_to_Product37_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out_to_Product37_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out_to_Subtract9_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out_to_Subtract9_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No20_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out_to_Subtract9_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out_to_Subtract9_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No21_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out_to_Subtract9_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out_to_Subtract9_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No22_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out_to_Subtract9_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out_to_Subtract9_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No23_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out_to_Subtract9_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out_to_Subtract9_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No249_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No24_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out_to_Product39_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out_to_Product39_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No3_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out_to_Subtract20_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out_to_Subtract20_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No30_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out_to_Subtract20_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out_to_Subtract20_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay3No206_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No31_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out_to_Subtract20_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out_to_Subtract20_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No32_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No254_out_to_Subtract20_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No255_out_to_Subtract20_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No33_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No256_out_to_Subtract20_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No257_out_to_Subtract20_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No34_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No258_out_to_Product220_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No259_out_to_Product220_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No260_out_to_Product220_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No261_out_to_Product220_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No262_out_to_Product220_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No263_out_to_Product220_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No264_out_to_Product323_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No265_out_to_Product323_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No266_out_to_Product323_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No267_out_to_Product323_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No268_out_to_Product323_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No269_out_to_Product323_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No270_out_to_Product323_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No271_out_to_Product323_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No272_out_to_Product325_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No273_out_to_Product325_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No274_out_to_Product325_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No275_out_to_Product325_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No276_out_to_Subtract26_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No277_out_to_Subtract26_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No278_out_to_Subtract26_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No279_out_to_Subtract26_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No280_out_to_Subtract26_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No281_out_to_Subtract26_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No282_out_to_Subtract26_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No283_out_to_Subtract26_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No284_out_to_Subtract26_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No285_out_to_Subtract26_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No286_out_to_Product55_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No287_out_to_Product55_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No288_out_to_Product55_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No289_out_to_Product55_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No290_out_to_Product55_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No291_out_to_Product55_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No292_out_to_Product226_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No293_out_to_Product226_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No294_out_to_Product226_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No295_out_to_Product226_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No296_out_to_Product326_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No297_out_to_Product326_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No298_out_to_Subtract29_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No299_out_to_Subtract29_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No300_out_to_Subtract29_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No301_out_to_Subtract29_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No302_out_to_Subtract29_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No303_out_to_Subtract29_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No304_out_to_Subtract29_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No305_out_to_Subtract29_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No306_out_to_Subtract29_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No307_out_to_Subtract29_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No308_out_to_Subtract33_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No309_out_to_Subtract33_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No310_out_to_Subtract33_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No311_out_to_Subtract33_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No312_out_to_Subtract33_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No313_out_to_Subtract33_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No314_out_to_Subtract33_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No315_out_to_Subtract33_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No316_out_to_Subtract33_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No317_out_to_Subtract33_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No318_out_to_Product237_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No319_out_to_Product237_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No320_out_to_Subtract38_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No321_out_to_Subtract38_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No322_out_to_Subtract38_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No323_out_to_Subtract38_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No324_out_to_Subtract38_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No325_out_to_Subtract38_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No326_out_to_Subtract38_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No327_out_to_Subtract38_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No328_out_to_Subtract38_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No329_out_to_Subtract38_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount141_instance: ModuloCounter_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount141_out);
x0_re_0_IEEE <= x0_re_0;
   x0_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_re_0_out,
                 X => x0_re_0_IEEE);
x0_im_0_IEEE <= x0_im_0;
   x0_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x0_im_0_out,
                 X => x0_im_0_IEEE);
x1_re_0_IEEE <= x1_re_0;
   x1_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_re_0_out,
                 X => x1_re_0_IEEE);
x1_im_0_IEEE <= x1_im_0;
   x1_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x1_im_0_out,
                 X => x1_im_0_IEEE);
x2_re_0_IEEE <= x2_re_0;
   x2_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_re_0_out,
                 X => x2_re_0_IEEE);
x2_im_0_IEEE <= x2_im_0;
   x2_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x2_im_0_out,
                 X => x2_im_0_IEEE);
x3_re_0_IEEE <= x3_re_0;
   x3_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_re_0_out,
                 X => x3_re_0_IEEE);
x3_im_0_IEEE <= x3_im_0;
   x3_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x3_im_0_out,
                 X => x3_im_0_IEEE);
x4_re_0_IEEE <= x4_re_0;
   x4_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_re_0_out,
                 X => x4_re_0_IEEE);
x4_im_0_IEEE <= x4_im_0;
   x4_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x4_im_0_out,
                 X => x4_im_0_IEEE);
x5_re_0_IEEE <= x5_re_0;
   x5_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_re_0_out,
                 X => x5_re_0_IEEE);
x5_im_0_IEEE <= x5_im_0;
   x5_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x5_im_0_out,
                 X => x5_im_0_IEEE);
x6_re_0_IEEE <= x6_re_0;
   x6_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_re_0_out,
                 X => x6_re_0_IEEE);
x6_im_0_IEEE <= x6_im_0;
   x6_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x6_im_0_out,
                 X => x6_im_0_IEEE);
x7_re_0_IEEE <= x7_re_0;
   x7_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_re_0_out,
                 X => x7_re_0_IEEE);
x7_im_0_IEEE <= x7_im_0;
   x7_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x7_im_0_out,
                 X => x7_im_0_IEEE);
x8_re_0_IEEE <= x8_re_0;
   x8_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_re_0_out,
                 X => x8_re_0_IEEE);
x8_im_0_IEEE <= x8_im_0;
   x8_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x8_im_0_out,
                 X => x8_im_0_IEEE);
x9_re_0_IEEE <= x9_re_0;
   x9_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_re_0_out,
                 X => x9_re_0_IEEE);
x9_im_0_IEEE <= x9_im_0;
   x9_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x9_im_0_out,
                 X => x9_im_0_IEEE);
x10_re_0_IEEE <= x10_re_0;
   x10_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_re_0_out,
                 X => x10_re_0_IEEE);
x10_im_0_IEEE <= x10_im_0;
   x10_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x10_im_0_out,
                 X => x10_im_0_IEEE);
x11_re_0_IEEE <= x11_re_0;
   x11_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_re_0_out,
                 X => x11_re_0_IEEE);
x11_im_0_IEEE <= x11_im_0;
   x11_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x11_im_0_out,
                 X => x11_im_0_IEEE);
x12_re_0_IEEE <= x12_re_0;
   x12_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_re_0_out,
                 X => x12_re_0_IEEE);
x12_im_0_IEEE <= x12_im_0;
   x12_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x12_im_0_out,
                 X => x12_im_0_IEEE);
x13_re_0_IEEE <= x13_re_0;
   x13_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_re_0_out,
                 X => x13_re_0_IEEE);
x13_im_0_IEEE <= x13_im_0;
   x13_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x13_im_0_out,
                 X => x13_im_0_IEEE);
x14_re_0_IEEE <= x14_re_0;
   x14_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_re_0_out,
                 X => x14_re_0_IEEE);
x14_im_0_IEEE <= x14_im_0;
   x14_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x14_im_0_out,
                 X => x14_im_0_IEEE);
x15_re_0_IEEE <= x15_re_0;
   x15_re_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_re_0_out,
                 X => x15_re_0_IEEE);
x15_im_0_IEEE <= x15_im_0;
   x15_im_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => x15_im_0_out,
                 X => x15_im_0_IEEE);
   y0_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_re_0_IEEE,
                 X => Delay1No_out);
y0_re_0 <= y0_re_0_IEEE;

SharedReg92_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg92_out;
SharedReg95_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg95_out;
SharedReg98_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg98_out;
SharedReg101_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg101_out;
SharedReg104_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg104_out;
   MUX_y0_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg92_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg95_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg98_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg101_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg104_out_to_MUX_y0_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y0_re_0_0_LUT_out,
                 oMux => MUX_y0_re_0_0_out);

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y0_re_0_0_out,
                 Y => Delay1No_out);
   y0_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y0_im_0_IEEE,
                 X => Delay1No1_out);
y0_im_0 <= y0_im_0_IEEE;

SharedReg107_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg107_out;
SharedReg112_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg112_out;
SharedReg117_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg117_out;
SharedReg122_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg122_out;
SharedReg127_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg127_out;
   MUX_y0_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg107_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg112_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg117_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg122_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg127_out_to_MUX_y0_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y0_im_0_0_LUT_out,
                 oMux => MUX_y0_im_0_0_out);

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y0_im_0_0_out,
                 Y => Delay1No1_out);
   y1_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_re_0_IEEE,
                 X => Delay1No2_out);
y1_re_0 <= y1_re_0_IEEE;

SharedReg132_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg132_out;
SharedReg137_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg137_out;
SharedReg142_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg142_out;
SharedReg147_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg147_out;
SharedReg152_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg152_out;
   MUX_y1_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg132_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg137_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg142_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg147_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg152_out_to_MUX_y1_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y1_re_0_0_LUT_out,
                 oMux => MUX_y1_re_0_0_out);

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y1_re_0_0_out,
                 Y => Delay1No2_out);
   y1_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y1_im_0_IEEE,
                 X => Delay1No3_out);
y1_im_0 <= y1_im_0_IEEE;

SharedReg32_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg32_out;
SharedReg38_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg38_out;
SharedReg44_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg44_out;
SharedReg50_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg50_out;
SharedReg56_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg56_out;
   MUX_y1_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg32_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg38_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg44_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg50_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg56_out_to_MUX_y1_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y1_im_0_0_LUT_out,
                 oMux => MUX_y1_im_0_0_out);

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y1_im_0_0_out,
                 Y => Delay1No3_out);
   y2_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_re_0_IEEE,
                 X => Delay1No4_out);
y2_re_0 <= y2_re_0_IEEE;

SharedReg62_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg62_out;
SharedReg68_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg68_out;
SharedReg74_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg74_out;
SharedReg80_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg80_out;
SharedReg86_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg86_out;
   MUX_y2_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg62_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg68_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg74_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg80_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg86_out_to_MUX_y2_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y2_re_0_0_LUT_out,
                 oMux => MUX_y2_re_0_0_out);

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y2_re_0_0_out,
                 Y => Delay1No4_out);
   y2_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y2_im_0_IEEE,
                 X => Delay1No5_out);
y2_im_0 <= y2_im_0_IEEE;

SharedReg92_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg92_out;
SharedReg95_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg95_out;
SharedReg98_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg98_out;
SharedReg101_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg101_out;
SharedReg104_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg104_out;
   MUX_y2_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg92_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg95_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg98_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg101_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg104_out_to_MUX_y2_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y2_im_0_0_LUT_out,
                 oMux => MUX_y2_im_0_0_out);

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y2_im_0_0_out,
                 Y => Delay1No5_out);
   y3_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_re_0_IEEE,
                 X => Delay1No6_out);
y3_re_0 <= y3_re_0_IEEE;

SharedReg92_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg92_out;
SharedReg95_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg95_out;
SharedReg98_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg98_out;
SharedReg101_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg101_out;
SharedReg104_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg104_out;
   MUX_y3_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg92_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg95_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg98_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg101_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg104_out_to_MUX_y3_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y3_re_0_0_LUT_out,
                 oMux => MUX_y3_re_0_0_out);

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y3_re_0_0_out,
                 Y => Delay1No6_out);
   y3_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y3_im_0_IEEE,
                 X => Delay1No7_out);
y3_im_0 <= y3_im_0_IEEE;

SharedReg107_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg107_out;
SharedReg112_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg112_out;
SharedReg117_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg117_out;
SharedReg122_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg122_out;
SharedReg127_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg127_out;
   MUX_y3_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg107_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg112_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg117_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg122_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg127_out_to_MUX_y3_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y3_im_0_0_LUT_out,
                 oMux => MUX_y3_im_0_0_out);

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y3_im_0_0_out,
                 Y => Delay1No7_out);
   y4_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_re_0_IEEE,
                 X => Delay1No8_out);
y4_re_0 <= y4_re_0_IEEE;

SharedReg132_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg132_out;
SharedReg137_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg137_out;
SharedReg142_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg142_out;
SharedReg147_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg147_out;
SharedReg152_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg152_out;
   MUX_y4_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg132_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg137_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg142_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg147_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg152_out_to_MUX_y4_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y4_re_0_0_LUT_out,
                 oMux => MUX_y4_re_0_0_out);

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y4_re_0_0_out,
                 Y => Delay1No8_out);
   y4_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y4_im_0_IEEE,
                 X => Delay1No9_out);
y4_im_0 <= y4_im_0_IEEE;

SharedReg157_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg157_out;
SharedReg165_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg165_out;
SharedReg173_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg173_out;
SharedReg181_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg181_out;
SharedReg189_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg189_out;
   MUX_y4_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg157_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg165_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg173_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg181_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg189_out_to_MUX_y4_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y4_im_0_0_LUT_out,
                 oMux => MUX_y4_im_0_0_out);

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y4_im_0_0_out,
                 Y => Delay1No9_out);
   y5_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_re_0_IEEE,
                 X => Delay1No10_out);
y5_re_0 <= y5_re_0_IEEE;

SharedReg62_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg62_out;
SharedReg68_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg68_out;
SharedReg74_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg74_out;
SharedReg80_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg80_out;
SharedReg86_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg86_out;
   MUX_y5_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg62_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg68_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg74_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg80_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg86_out_to_MUX_y5_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y5_re_0_0_LUT_out,
                 oMux => MUX_y5_re_0_0_out);

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y5_re_0_0_out,
                 Y => Delay1No10_out);
   y5_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y5_im_0_IEEE,
                 X => Delay1No11_out);
y5_im_0 <= y5_im_0_IEEE;

SharedReg92_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg92_out;
SharedReg95_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg95_out;
SharedReg98_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg98_out;
SharedReg101_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg101_out;
SharedReg104_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg104_out;
   MUX_y5_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg92_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg95_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg98_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg101_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg104_out_to_MUX_y5_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y5_im_0_0_LUT_out,
                 oMux => MUX_y5_im_0_0_out);

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y5_im_0_0_out,
                 Y => Delay1No11_out);
   y6_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_re_0_IEEE,
                 X => Delay1No12_out);
y6_re_0 <= y6_re_0_IEEE;

SharedReg107_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg107_out;
SharedReg112_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg112_out;
SharedReg117_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg117_out;
SharedReg122_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg122_out;
SharedReg127_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg127_out;
   MUX_y6_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg107_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg112_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg117_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg122_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg127_out_to_MUX_y6_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y6_re_0_0_LUT_out,
                 oMux => MUX_y6_re_0_0_out);

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y6_re_0_0_out,
                 Y => Delay1No12_out);
   y6_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y6_im_0_IEEE,
                 X => Delay1No13_out);
y6_im_0 <= y6_im_0_IEEE;

SharedReg132_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg132_out;
SharedReg137_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg137_out;
SharedReg142_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg142_out;
SharedReg147_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg147_out;
SharedReg152_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg152_out;
   MUX_y6_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg132_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg137_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg142_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg147_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg152_out_to_MUX_y6_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y6_im_0_0_LUT_out,
                 oMux => MUX_y6_im_0_0_out);

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y6_im_0_0_out,
                 Y => Delay1No13_out);
   y7_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_re_0_IEEE,
                 X => Delay1No14_out);
y7_re_0 <= y7_re_0_IEEE;

SharedReg107_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg107_out;
SharedReg112_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg112_out;
SharedReg117_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg117_out;
SharedReg122_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg122_out;
SharedReg127_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg127_out;
   MUX_y7_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg107_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg112_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg117_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg122_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg127_out_to_MUX_y7_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y7_re_0_0_LUT_out,
                 oMux => MUX_y7_re_0_0_out);

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y7_re_0_0_out,
                 Y => Delay1No14_out);
   y7_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y7_im_0_IEEE,
                 X => Delay1No15_out);
y7_im_0 <= y7_im_0_IEEE;

SharedReg132_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg132_out;
SharedReg137_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg137_out;
SharedReg142_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg142_out;
SharedReg147_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg147_out;
SharedReg152_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg152_out;
   MUX_y7_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg132_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg137_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg142_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg147_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg152_out_to_MUX_y7_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y7_im_0_0_LUT_out,
                 oMux => MUX_y7_im_0_0_out);

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y7_im_0_0_out,
                 Y => Delay1No15_out);
   y8_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_re_0_IEEE,
                 X => Delay1No16_out);
y8_re_0 <= y8_re_0_IEEE;

SharedReg704_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg704_out;
SharedReg710_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg710_out;
SharedReg716_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg716_out;
SharedReg722_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg722_out;
SharedReg728_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg728_out;
   MUX_y8_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg704_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg710_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg716_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg722_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg728_out_to_MUX_y8_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y8_re_0_0_LUT_out,
                 oMux => MUX_y8_re_0_0_out);

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y8_re_0_0_out,
                 Y => Delay1No16_out);
   y8_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y8_im_0_IEEE,
                 X => Delay1No17_out);
y8_im_0 <= y8_im_0_IEEE;

SharedReg736_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg736_out;
SharedReg744_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg744_out;
SharedReg752_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg752_out;
SharedReg760_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg760_out;
SharedReg768_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg768_out;
   MUX_y8_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg736_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg744_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg752_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg760_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg768_out_to_MUX_y8_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y8_im_0_0_LUT_out,
                 oMux => MUX_y8_im_0_0_out);

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y8_im_0_0_out,
                 Y => Delay1No17_out);
   y9_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_re_0_IEEE,
                 X => Delay1No18_out);
y9_re_0 <= y9_re_0_IEEE;

SharedReg704_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg704_out;
SharedReg710_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg710_out;
SharedReg716_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg716_out;
SharedReg722_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg722_out;
SharedReg728_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg728_out;
   MUX_y9_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg704_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg710_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg716_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg722_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg728_out_to_MUX_y9_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y9_re_0_0_LUT_out,
                 oMux => MUX_y9_re_0_0_out);

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y9_re_0_0_out,
                 Y => Delay1No18_out);
   y9_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y9_im_0_IEEE,
                 X => Delay1No19_out);
y9_im_0 <= y9_im_0_IEEE;

SharedReg736_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg736_out;
SharedReg744_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg744_out;
SharedReg752_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg752_out;
SharedReg760_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg760_out;
SharedReg768_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg768_out;
   MUX_y9_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg736_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg744_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg752_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg760_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg768_out_to_MUX_y9_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y9_im_0_0_LUT_out,
                 oMux => MUX_y9_im_0_0_out);

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y9_im_0_0_out,
                 Y => Delay1No19_out);
   y10_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_re_0_IEEE,
                 X => Delay1No20_out);
y10_re_0 <= y10_re_0_IEEE;

SharedReg574_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg574_out;
SharedReg579_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg579_out;
SharedReg584_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg584_out;
SharedReg589_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg589_out;
SharedReg594_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg594_out;
   MUX_y10_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg574_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg579_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg584_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg589_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg594_out_to_MUX_y10_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y10_re_0_0_LUT_out,
                 oMux => MUX_y10_re_0_0_out);

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y10_re_0_0_out,
                 Y => Delay1No20_out);
   y10_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y10_im_0_IEEE,
                 X => Delay1No21_out);
y10_im_0 <= y10_im_0_IEEE;

SharedReg637_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg637_out;
SharedReg642_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg642_out;
SharedReg647_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg647_out;
SharedReg652_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg652_out;
SharedReg657_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg657_out;
   MUX_y10_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg637_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg642_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg647_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg652_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg657_out_to_MUX_y10_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y10_im_0_0_LUT_out,
                 oMux => MUX_y10_im_0_0_out);

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y10_im_0_0_out,
                 Y => Delay1No21_out);
   y11_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_re_0_IEEE,
                 X => Delay1No22_out);
y11_re_0 <= y11_re_0_IEEE;

SharedReg704_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg704_out;
SharedReg710_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg710_out;
SharedReg716_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg716_out;
SharedReg722_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg722_out;
SharedReg728_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg728_out;
   MUX_y11_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg704_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg710_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg716_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg722_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg728_out_to_MUX_y11_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y11_re_0_0_LUT_out,
                 oMux => MUX_y11_re_0_0_out);

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y11_re_0_0_out,
                 Y => Delay1No22_out);
   y11_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y11_im_0_IEEE,
                 X => Delay1No23_out);
y11_im_0 <= y11_im_0_IEEE;

SharedReg736_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg736_out;
SharedReg744_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg744_out;
SharedReg752_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg752_out;
SharedReg760_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg760_out;
SharedReg768_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg768_out;
   MUX_y11_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg736_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg744_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg752_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg760_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg768_out_to_MUX_y11_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y11_im_0_0_LUT_out,
                 oMux => MUX_y11_im_0_0_out);

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y11_im_0_0_out,
                 Y => Delay1No23_out);
   y12_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_re_0_IEEE,
                 X => Delay1No24_out);
y12_re_0 <= y12_re_0_IEEE;

SharedReg736_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg736_out;
SharedReg744_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg744_out;
SharedReg752_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg752_out;
SharedReg760_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg760_out;
SharedReg768_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg768_out;
   MUX_y12_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg736_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg744_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg752_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg760_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg768_out_to_MUX_y12_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y12_re_0_0_LUT_out,
                 oMux => MUX_y12_re_0_0_out);

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y12_re_0_0_out,
                 Y => Delay1No24_out);
   y12_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y12_im_0_IEEE,
                 X => Delay1No25_out);
y12_im_0 <= y12_im_0_IEEE;

SharedReg546_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg546_out;
SharedReg551_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg551_out;
SharedReg556_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg556_out;
SharedReg561_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg566_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg566_out;
   MUX_y12_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg546_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg551_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg556_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg566_out_to_MUX_y12_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y12_im_0_0_LUT_out,
                 oMux => MUX_y12_im_0_0_out);

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y12_im_0_0_out,
                 Y => Delay1No25_out);
   y13_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_re_0_IEEE,
                 X => Delay1No26_out);
y13_re_0 <= y13_re_0_IEEE;

SharedReg637_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg637_out;
SharedReg642_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg642_out;
SharedReg647_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg647_out;
SharedReg652_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg652_out;
SharedReg657_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg657_out;
   MUX_y13_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg637_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg642_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg647_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg652_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg657_out_to_MUX_y13_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y13_re_0_0_LUT_out,
                 oMux => MUX_y13_re_0_0_out);

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y13_re_0_0_out,
                 Y => Delay1No26_out);
   y13_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y13_im_0_IEEE,
                 X => Delay1No27_out);
y13_im_0 <= y13_im_0_IEEE;

SharedReg679_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg679_out;
SharedReg684_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg684_out;
SharedReg689_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg689_out;
SharedReg694_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg694_out;
SharedReg699_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg699_out;
   MUX_y13_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg679_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg684_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg689_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg694_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg699_out_to_MUX_y13_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y13_im_0_0_LUT_out,
                 oMux => MUX_y13_im_0_0_out);

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y13_im_0_0_out,
                 Y => Delay1No27_out);
   y14_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_re_0_IEEE,
                 X => Delay1No28_out);
y14_re_0 <= y14_re_0_IEEE;

SharedReg679_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg679_out;
SharedReg684_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg684_out;
SharedReg689_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg689_out;
SharedReg694_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg694_out;
SharedReg699_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg699_out;
   MUX_y14_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg679_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg684_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg689_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg694_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg699_out_to_MUX_y14_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y14_re_0_0_LUT_out,
                 oMux => MUX_y14_re_0_0_out);

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y14_re_0_0_out,
                 Y => Delay1No28_out);
   y14_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y14_im_0_IEEE,
                 X => Delay1No29_out);
y14_im_0 <= y14_im_0_IEEE;

SharedReg704_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg704_out;
SharedReg710_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg710_out;
SharedReg716_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg716_out;
SharedReg722_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg722_out;
SharedReg728_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg728_out;
   MUX_y14_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg704_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg710_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg716_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg722_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg728_out_to_MUX_y14_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y14_im_0_0_LUT_out,
                 oMux => MUX_y14_im_0_0_out);

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y14_im_0_0_out,
                 Y => Delay1No29_out);
   y15_re_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_re_0_IEEE,
                 X => Delay1No30_out);
y15_re_0 <= y15_re_0_IEEE;

SharedReg704_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast <= SharedReg704_out;
SharedReg710_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast <= SharedReg710_out;
SharedReg716_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast <= SharedReg716_out;
SharedReg722_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast <= SharedReg722_out;
SharedReg728_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast <= SharedReg728_out;
   MUX_y15_re_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg704_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg710_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg716_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg722_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg728_out_to_MUX_y15_re_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y15_re_0_0_LUT_out,
                 oMux => MUX_y15_re_0_0_out);

   Delay1No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y15_re_0_0_out,
                 Y => Delay1No30_out);
   y15_im_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => y15_im_0_IEEE,
                 X => Delay1No31_out);
y15_im_0 <= y15_im_0_IEEE;

SharedReg736_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast <= SharedReg736_out;
SharedReg744_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast <= SharedReg744_out;
SharedReg752_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast <= SharedReg752_out;
SharedReg760_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast <= SharedReg760_out;
SharedReg768_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast <= SharedReg768_out;
   MUX_y15_im_0_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg736_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg744_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg752_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg760_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg768_out_to_MUX_y15_im_0_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_y15_im_0_0_LUT_out,
                 oMux => MUX_y15_im_0_0_out);

   Delay1No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_y15_im_0_0_out,
                 Y => Delay1No31_out);

Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast <= Delay1No32_out;
Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast <= Delay1No33_out;
   Add2_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_0_impl_out,
                 X => Delay1No32_out_to_Add2_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No33_out_to_Add2_0_impl_parent_implementedSystem_port_1_cast);

SharedReg201_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg201_out;
SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg12_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg12_out;
SharedReg576_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg576_out;
SharedReg546_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg546_out;
SharedReg327_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg327_out;
SharedReg306_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg306_out;
SharedReg135_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg135_out;
SharedReg546_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg546_out;
SharedReg330_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg330_out;
SharedReg160_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg160_out;
SharedReg162_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg162_out;
SharedReg326_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg326_out;
SharedReg198_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg198_out;
   MUX_Add2_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg201_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg160_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg162_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg326_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg198_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg12_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg576_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg546_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg327_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg306_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg135_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg546_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg330_out_to_MUX_Add2_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add2_0_impl_0_out);

   Delay1No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_0_impl_0_out,
                 Y => Delay1No32_out);

SharedReg133_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg133_out;
SharedReg16_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg28_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg28_out;
SharedReg490_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg490_out;
SharedReg574_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg574_out;
SharedReg546_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg546_out;
SharedReg305_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg305_out;
SharedReg161_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg161_out;
SharedReg574_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg574_out;
SharedReg546_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg546_out;
SharedReg132_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg132_out;
SharedReg32_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg32_out;
SharedReg491_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg491_out;
SharedReg200_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg200_out;
   MUX_Add2_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg133_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg132_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg32_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg491_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg200_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg28_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg490_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg574_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg546_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg305_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg161_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg574_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg546_out_to_MUX_Add2_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add2_0_impl_1_out);

   Delay1No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_0_impl_1_out,
                 Y => Delay1No33_out);

Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast <= Delay1No34_out;
Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast <= Delay1No35_out;
   Add2_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_1_impl_out,
                 X => Delay1No34_out_to_Add2_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No35_out_to_Add2_1_impl_parent_implementedSystem_port_1_cast);

SharedReg170_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg170_out;
SharedReg333_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg333_out;
SharedReg206_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg206_out;
SharedReg209_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg209_out;
SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg_out;
SharedReg12_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg12_out;
SharedReg581_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg581_out;
SharedReg551_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg551_out;
SharedReg334_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg334_out;
SharedReg320_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg320_out;
SharedReg140_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg140_out;
SharedReg551_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg551_out;
SharedReg337_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg337_out;
SharedReg168_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg168_out;
   MUX_Add2_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg170_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg333_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg140_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg551_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg337_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg168_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg206_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg209_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg12_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg581_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg551_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg334_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg320_out_to_MUX_Add2_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add2_1_impl_0_out);

   Delay1No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_1_impl_0_out,
                 Y => Delay1No34_out);

SharedReg38_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg38_out;
SharedReg498_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg498_out;
SharedReg208_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg208_out;
SharedReg138_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg138_out;
SharedReg16_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg16_out;
SharedReg28_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg28_out;
SharedReg497_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg497_out;
SharedReg579_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg579_out;
SharedReg551_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg551_out;
SharedReg319_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg319_out;
SharedReg169_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg169_out;
SharedReg579_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg579_out;
SharedReg551_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg551_out;
SharedReg137_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg137_out;
   MUX_Add2_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg38_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg498_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg169_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg579_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg551_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg137_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg208_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg138_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg16_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg28_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg497_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg579_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg551_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg319_out_to_MUX_Add2_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add2_1_impl_1_out);

   Delay1No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_1_impl_1_out,
                 Y => Delay1No35_out);

Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast <= Delay1No36_out;
Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast <= Delay1No37_out;
   Add2_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_2_impl_out,
                 X => Delay1No36_out_to_Add2_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No37_out_to_Add2_2_impl_parent_implementedSystem_port_1_cast);

SharedReg556_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg556_out;
SharedReg344_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg344_out;
SharedReg176_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg176_out;
SharedReg178_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg178_out;
SharedReg340_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg340_out;
SharedReg214_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg214_out;
SharedReg217_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg217_out;
SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg_out;
SharedReg12_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg12_out;
SharedReg586_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg586_out;
SharedReg556_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg556_out;
SharedReg341_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg341_out;
SharedReg311_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg311_out;
SharedReg145_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg145_out;
   MUX_Add2_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg556_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg344_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg556_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg341_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg311_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg145_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg176_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg178_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg340_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg214_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg217_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg12_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg586_out_to_MUX_Add2_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add2_2_impl_0_out);

   Delay1No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_2_impl_0_out,
                 Y => Delay1No36_out);

SharedReg584_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg584_out;
SharedReg556_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg556_out;
SharedReg142_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg142_out;
SharedReg44_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg44_out;
SharedReg505_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg505_out;
SharedReg216_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg216_out;
SharedReg143_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg143_out;
SharedReg16_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg16_out;
SharedReg28_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg28_out;
SharedReg504_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg504_out;
SharedReg584_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg584_out;
SharedReg556_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg556_out;
SharedReg369_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg369_out;
SharedReg177_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg177_out;
   MUX_Add2_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg584_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg556_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg584_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg556_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg369_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg177_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg142_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg44_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg505_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg216_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg143_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg16_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg28_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg504_out_to_MUX_Add2_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add2_2_impl_1_out);

   Delay1No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_2_impl_1_out,
                 Y => Delay1No37_out);

Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast <= Delay1No38_out;
Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast <= Delay1No39_out;
   Add2_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_3_impl_out,
                 X => Delay1No38_out_to_Add2_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No39_out_to_Add2_3_impl_parent_implementedSystem_port_1_cast);

SharedReg348_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg348_out;
SharedReg316_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg316_out;
SharedReg150_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg150_out;
SharedReg561_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg351_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg351_out;
SharedReg184_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg184_out;
SharedReg186_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg186_out;
SharedReg347_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg347_out;
SharedReg222_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg222_out;
SharedReg225_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg225_out;
SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg_out;
SharedReg12_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg12_out;
SharedReg591_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg591_out;
SharedReg561_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg561_out;
   MUX_Add2_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg348_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg316_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg12_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg591_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg561_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg150_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg351_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg184_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg186_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg347_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg222_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg225_out_to_MUX_Add2_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add2_3_impl_0_out);

   Delay1No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_3_impl_0_out,
                 Y => Delay1No38_out);

SharedReg561_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg372_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg372_out;
SharedReg185_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg185_out;
SharedReg589_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg589_out;
SharedReg561_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg561_out;
SharedReg147_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg147_out;
SharedReg50_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg50_out;
SharedReg512_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg512_out;
SharedReg224_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg224_out;
SharedReg148_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg148_out;
SharedReg16_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg16_out;
SharedReg28_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg28_out;
SharedReg511_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg511_out;
SharedReg589_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg589_out;
   MUX_Add2_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg372_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg16_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg28_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg511_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg589_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg185_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg589_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg561_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg147_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg50_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg512_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg224_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg148_out_to_MUX_Add2_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add2_3_impl_1_out);

   Delay1No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_3_impl_1_out,
                 Y => Delay1No39_out);

Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast <= Delay1No40_out;
Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast <= Delay1No41_out;
   Add2_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add2_4_impl_out,
                 X => Delay1No40_out_to_Add2_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No41_out_to_Add2_4_impl_parent_implementedSystem_port_1_cast);

SharedReg596_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg596_out;
SharedReg566_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg566_out;
SharedReg355_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg355_out;
SharedReg325_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg325_out;
SharedReg155_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg155_out;
SharedReg566_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg566_out;
SharedReg358_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg358_out;
SharedReg192_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg192_out;
SharedReg194_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg194_out;
SharedReg354_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg354_out;
SharedReg230_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg230_out;
SharedReg233_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg233_out;
SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg_out;
SharedReg12_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg12_out;
   MUX_Add2_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg596_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg566_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg230_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg233_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg12_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg355_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg325_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg155_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg566_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg358_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg192_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg194_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg354_out_to_MUX_Add2_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add2_4_impl_0_out);

   Delay1No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_4_impl_0_out,
                 Y => Delay1No40_out);

SharedReg518_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg518_out;
SharedReg594_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg594_out;
SharedReg566_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg566_out;
SharedReg302_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg302_out;
SharedReg193_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg193_out;
SharedReg594_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg594_out;
SharedReg566_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg566_out;
SharedReg152_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg152_out;
SharedReg56_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg56_out;
SharedReg519_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg519_out;
SharedReg232_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg232_out;
SharedReg153_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg153_out;
SharedReg16_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg16_out;
SharedReg28_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg28_out;
   MUX_Add2_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg518_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg594_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg232_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg153_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg16_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg28_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg566_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg302_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg193_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg594_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg566_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg152_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg56_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg519_out_to_MUX_Add2_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add2_4_impl_1_out);

   Delay1No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add2_4_impl_1_out,
                 Y => Delay1No41_out);

Delay1No42_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast <= Delay1No42_out;
Delay1No43_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast <= Delay1No43_out;
   Add11_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_0_impl_out,
                 X => Delay1No42_out_to_Add11_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No43_out_to_Add11_0_impl_parent_implementedSystem_port_1_cast);

SharedReg492_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg492_out;
SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg6_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg6_out;
SharedReg198_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg198_out;
SharedReg197_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg197_out;
SharedReg158_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg158_out;
SharedReg376_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg376_out;
SharedReg550_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg550_out;
SharedReg326_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg326_out;
SharedReg332_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg332_out;
SharedReg494_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg494_out;
SharedReg203_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg203_out;
SharedReg107_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg107_out;
SharedReg490_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg490_out;
   MUX_Add11_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg492_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg494_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg203_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg107_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg490_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg6_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg198_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg197_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg158_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg376_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg550_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg326_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg332_out_to_MUX_Add11_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add11_0_impl_0_out);

   Delay1No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_0_impl_0_out,
                 Y => Delay1No42_out);

SharedReg326_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg326_out;
SharedReg17_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg17_out;
SharedReg22_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg22_out;
SharedReg197_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg197_out;
SharedReg237_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg237_out;
SharedReg197_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg197_out;
SharedReg393_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg393_out;
SharedReg496_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg496_out;
SharedReg490_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg490_out;
SharedReg331_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg331_out;
SharedReg326_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg326_out;
SharedReg237_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg237_out;
SharedReg63_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg63_out;
SharedReg549_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg549_out;
   MUX_Add11_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg326_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg17_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg326_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg237_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg63_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg549_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg22_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg197_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg237_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg197_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg393_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg496_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg490_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg331_out_to_MUX_Add11_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add11_0_impl_1_out);

   Delay1No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_0_impl_1_out,
                 Y => Delay1No43_out);

Delay1No44_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast <= Delay1No44_out;
Delay1No45_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast <= Delay1No45_out;
   Add11_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_1_impl_out,
                 X => Delay1No44_out_to_Add11_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No45_out_to_Add11_1_impl_parent_implementedSystem_port_1_cast);

SharedReg211_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg211_out;
SharedReg112_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg112_out;
SharedReg497_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg497_out;
SharedReg499_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg499_out;
SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1_out;
SharedReg6_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg6_out;
SharedReg206_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg206_out;
SharedReg205_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg205_out;
SharedReg166_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg166_out;
SharedReg364_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg364_out;
SharedReg555_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg555_out;
SharedReg333_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg333_out;
SharedReg339_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg339_out;
SharedReg501_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg501_out;
   MUX_Add11_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg211_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg112_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg555_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg333_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg339_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg501_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg497_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg499_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg6_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg206_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg205_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg166_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg364_out_to_MUX_Add11_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add11_1_impl_0_out);

   Delay1No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_1_impl_0_out,
                 Y => Delay1No44_out);

SharedReg246_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg246_out;
SharedReg69_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg69_out;
SharedReg554_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg554_out;
SharedReg333_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg333_out;
SharedReg17_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg17_out;
SharedReg22_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg22_out;
SharedReg205_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg205_out;
SharedReg246_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg246_out;
SharedReg205_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg205_out;
SharedReg379_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg379_out;
SharedReg503_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg503_out;
SharedReg497_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg497_out;
SharedReg338_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg338_out;
SharedReg333_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg333_out;
   MUX_Add11_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg246_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg69_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg503_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg497_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg338_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg333_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg554_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg333_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg17_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg22_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg205_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg246_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg205_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg379_out_to_MUX_Add11_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add11_1_impl_1_out);

   Delay1No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_1_impl_1_out,
                 Y => Delay1No45_out);

Delay1No46_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast <= Delay1No46_out;
Delay1No47_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast <= Delay1No47_out;
   Add11_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_2_impl_out,
                 X => Delay1No46_out_to_Add11_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No47_out_to_Add11_2_impl_parent_implementedSystem_port_1_cast);

SharedReg340_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg340_out;
SharedReg346_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg346_out;
SharedReg508_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg508_out;
SharedReg219_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg219_out;
SharedReg117_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg117_out;
SharedReg504_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg504_out;
SharedReg506_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg506_out;
SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1_out;
SharedReg6_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg6_out;
SharedReg214_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg214_out;
SharedReg213_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg213_out;
SharedReg174_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg174_out;
SharedReg382_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg382_out;
SharedReg560_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg560_out;
   MUX_Add11_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg340_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg346_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg213_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg174_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg382_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg560_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg508_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg219_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg117_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg504_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg506_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg6_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg214_out_to_MUX_Add11_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add11_2_impl_0_out);

   Delay1No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_2_impl_0_out,
                 Y => Delay1No46_out);

SharedReg504_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg504_out;
SharedReg345_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg345_out;
SharedReg340_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg340_out;
SharedReg255_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg255_out;
SharedReg75_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg75_out;
SharedReg559_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg559_out;
SharedReg340_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg340_out;
SharedReg17_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg17_out;
SharedReg22_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg22_out;
SharedReg213_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg213_out;
SharedReg255_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg255_out;
SharedReg213_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg213_out;
SharedReg400_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg400_out;
SharedReg510_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg510_out;
   MUX_Add11_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg504_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg345_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg255_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg213_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg400_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg510_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg340_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg255_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg75_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg559_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg340_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg17_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg22_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg213_out_to_MUX_Add11_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add11_2_impl_1_out);

   Delay1No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_2_impl_1_out,
                 Y => Delay1No47_out);

Delay1No48_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast <= Delay1No48_out;
Delay1No49_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast <= Delay1No49_out;
   Add11_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_3_impl_out,
                 X => Delay1No48_out_to_Add11_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No49_out_to_Add11_3_impl_parent_implementedSystem_port_1_cast);

SharedReg182_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg182_out;
SharedReg370_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg370_out;
SharedReg565_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg565_out;
SharedReg347_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg347_out;
SharedReg353_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg353_out;
SharedReg515_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg515_out;
SharedReg227_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg227_out;
SharedReg122_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg122_out;
SharedReg511_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg511_out;
SharedReg513_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg513_out;
SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1_out;
SharedReg6_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg6_out;
SharedReg222_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg222_out;
SharedReg221_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg221_out;
   MUX_Add11_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg182_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg370_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg6_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg222_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg221_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg565_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg347_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg353_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg515_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg227_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg122_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg511_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg513_out_to_MUX_Add11_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add11_3_impl_0_out);

   Delay1No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_3_impl_0_out,
                 Y => Delay1No48_out);

SharedReg221_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg221_out;
SharedReg386_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg386_out;
SharedReg517_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg517_out;
SharedReg511_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg511_out;
SharedReg352_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg352_out;
SharedReg347_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg347_out;
SharedReg264_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg264_out;
SharedReg81_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg81_out;
SharedReg564_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg564_out;
SharedReg347_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg347_out;
SharedReg17_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg17_out;
SharedReg22_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg22_out;
SharedReg221_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg221_out;
SharedReg264_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg264_out;
   MUX_Add11_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg221_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg386_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg17_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg22_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg221_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg264_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg517_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg511_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg352_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg347_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg264_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg81_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg564_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg347_out_to_MUX_Add11_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add11_3_impl_1_out);

   Delay1No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_3_impl_1_out,
                 Y => Delay1No49_out);

Delay1No50_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast <= Delay1No50_out;
Delay1No51_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast <= Delay1No51_out;
   Add11_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add11_4_impl_out,
                 X => Delay1No50_out_to_Add11_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No51_out_to_Add11_4_impl_parent_implementedSystem_port_1_cast);

SharedReg230_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg230_out;
SharedReg229_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg229_out;
SharedReg190_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg190_out;
SharedReg390_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg390_out;
SharedReg570_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg570_out;
SharedReg354_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg354_out;
SharedReg360_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg360_out;
SharedReg522_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg522_out;
SharedReg235_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg235_out;
SharedReg127_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg127_out;
SharedReg518_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg518_out;
SharedReg520_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg520_out;
SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1_out;
SharedReg6_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg6_out;
   MUX_Add11_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg230_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg229_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg518_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg520_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg6_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg190_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg390_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg570_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg354_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg360_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg522_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg235_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg127_out_to_MUX_Add11_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add11_4_impl_0_out);

   Delay1No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_4_impl_0_out,
                 Y => Delay1No50_out);

SharedReg229_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg229_out;
SharedReg273_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg273_out;
SharedReg229_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg229_out;
SharedReg407_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg407_out;
SharedReg524_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg524_out;
SharedReg518_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg518_out;
SharedReg359_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg359_out;
SharedReg354_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg354_out;
SharedReg273_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg273_out;
SharedReg87_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg87_out;
SharedReg569_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg569_out;
SharedReg354_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg354_out;
SharedReg17_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg17_out;
SharedReg22_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg22_out;
   MUX_Add11_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg229_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg273_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg569_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg354_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg17_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg22_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg229_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg407_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg524_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg518_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg359_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg354_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg273_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg87_out_to_MUX_Add11_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add11_4_impl_1_out);

   Delay1No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add11_4_impl_1_out,
                 Y => Delay1No51_out);

Delay1No52_out_to_Add3_0_impl_parent_implementedSystem_port_0_cast <= Delay1No52_out;
Delay1No53_out_to_Add3_0_impl_parent_implementedSystem_port_1_cast <= Delay1No53_out;
   Add3_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_0_impl_out,
                 X => Delay1No52_out_to_Add3_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No53_out_to_Add3_0_impl_parent_implementedSystem_port_1_cast);

SharedReg547_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg547_out;
SharedReg2_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg2_out;
SharedReg7_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg7_out;
SharedReg305_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg305_out;
SharedReg548_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg548_out;
SharedReg328_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg328_out;
SharedReg434_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg434_out;
SharedReg202_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg202_out;
SharedReg92_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg92_out;
SharedReg495_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg495_out;
SharedReg158_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg158_out;
SharedReg495_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg495_out;
SharedReg547_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg547_out;
SharedReg238_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg238_out;
   MUX_Add3_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg547_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg2_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg158_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg495_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg547_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg238_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg7_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg305_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg548_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg328_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg434_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg202_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg92_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg495_out_to_MUX_Add3_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add3_0_impl_0_out);

   Delay1No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_0_impl_0_out,
                 Y => Delay1No52_out);

SharedReg641_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg641_out;
SharedReg18_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg23_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg23_out;
SharedReg433_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg433_out;
SharedReg490_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg490_out;
SharedReg574_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg574_out;
SharedReg395_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg395_out;
SharedReg136_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg136_out;
SharedReg107_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg107_out;
SharedReg683_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg683_out;
SharedReg157_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg157_out;
SharedReg326_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg326_out;
SharedReg638_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg638_out;
SharedReg240_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg240_out;
   MUX_Add3_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg641_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg157_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg326_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg638_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg240_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg23_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg433_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg490_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg574_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg395_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg136_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg107_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg683_out_to_MUX_Add3_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add3_0_impl_1_out);

   Delay1No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_0_impl_1_out,
                 Y => Delay1No53_out);

Delay1No54_out_to_Add3_1_impl_parent_implementedSystem_port_0_cast <= Delay1No54_out;
Delay1No55_out_to_Add3_1_impl_parent_implementedSystem_port_1_cast <= Delay1No55_out;
   Add3_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_1_impl_out,
                 X => Delay1No54_out_to_Add3_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No55_out_to_Add3_1_impl_parent_implementedSystem_port_1_cast);

SharedReg502_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg502_out;
SharedReg552_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg552_out;
SharedReg247_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg247_out;
SharedReg552_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg552_out;
SharedReg2_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg2_out;
SharedReg7_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg7_out;
SharedReg319_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg319_out;
SharedReg553_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg553_out;
SharedReg335_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg335_out;
SharedReg438_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg438_out;
SharedReg210_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg210_out;
SharedReg95_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg95_out;
SharedReg502_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg502_out;
SharedReg166_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg166_out;
   MUX_Add3_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg502_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg552_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg210_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg95_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg502_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg166_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg247_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg552_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg2_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg7_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg319_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg553_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg335_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg438_out_to_MUX_Add3_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add3_1_impl_0_out);

   Delay1No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_1_impl_0_out,
                 Y => Delay1No54_out);

SharedReg333_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg333_out;
SharedReg643_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg643_out;
SharedReg249_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg249_out;
SharedReg646_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg646_out;
SharedReg18_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg18_out;
SharedReg23_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg23_out;
SharedReg417_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg417_out;
SharedReg497_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg497_out;
SharedReg579_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg579_out;
SharedReg398_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg398_out;
SharedReg141_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg141_out;
SharedReg112_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg112_out;
SharedReg688_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg688_out;
SharedReg165_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg165_out;
   MUX_Add3_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg333_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg643_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg141_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg112_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg688_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg165_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg249_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg646_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg18_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg23_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg417_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg497_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg579_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg398_out_to_MUX_Add3_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add3_1_impl_1_out);

   Delay1No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_1_impl_1_out,
                 Y => Delay1No55_out);

Delay1No56_out_to_Add3_2_impl_parent_implementedSystem_port_0_cast <= Delay1No56_out;
Delay1No57_out_to_Add3_2_impl_parent_implementedSystem_port_1_cast <= Delay1No57_out;
   Add3_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_2_impl_out,
                 X => Delay1No56_out_to_Add3_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No57_out_to_Add3_2_impl_parent_implementedSystem_port_1_cast);

SharedReg98_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg98_out;
SharedReg509_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg509_out;
SharedReg174_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg174_out;
SharedReg509_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg509_out;
SharedReg557_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg557_out;
SharedReg256_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg256_out;
SharedReg557_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg557_out;
SharedReg2_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg2_out;
SharedReg7_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg7_out;
SharedReg369_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg369_out;
SharedReg558_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg558_out;
SharedReg342_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg342_out;
SharedReg460_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg460_out;
SharedReg218_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg218_out;
   MUX_Add3_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg98_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg509_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg558_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg342_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg460_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg218_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg174_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg509_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg557_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg256_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg557_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg2_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg7_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg369_out_to_MUX_Add3_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add3_2_impl_0_out);

   Delay1No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_2_impl_0_out,
                 Y => Delay1No56_out);

SharedReg117_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg117_out;
SharedReg693_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg693_out;
SharedReg173_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg173_out;
SharedReg340_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg340_out;
SharedReg648_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg648_out;
SharedReg258_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg258_out;
SharedReg651_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg651_out;
SharedReg18_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg18_out;
SharedReg23_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg23_out;
SharedReg442_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg442_out;
SharedReg504_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg504_out;
SharedReg584_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg584_out;
SharedReg420_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg420_out;
SharedReg146_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg146_out;
   MUX_Add3_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg117_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg693_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg504_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg584_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg420_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg146_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg173_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg340_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg648_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg258_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg651_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg18_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg23_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg442_out_to_MUX_Add3_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add3_2_impl_1_out);

   Delay1No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_2_impl_1_out,
                 Y => Delay1No57_out);

Delay1No58_out_to_Add3_3_impl_parent_implementedSystem_port_0_cast <= Delay1No58_out;
Delay1No59_out_to_Add3_3_impl_parent_implementedSystem_port_1_cast <= Delay1No59_out;
   Add3_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_3_impl_out,
                 X => Delay1No58_out_to_Add3_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No59_out_to_Add3_3_impl_parent_implementedSystem_port_1_cast);

SharedReg349_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg349_out;
SharedReg465_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg465_out;
SharedReg226_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg226_out;
SharedReg101_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg101_out;
SharedReg516_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg516_out;
SharedReg182_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg182_out;
SharedReg516_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg516_out;
SharedReg562_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg562_out;
SharedReg265_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg265_out;
SharedReg562_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg562_out;
SharedReg2_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg2_out;
SharedReg7_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg7_out;
SharedReg372_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg372_out;
SharedReg563_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg563_out;
   MUX_Add3_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg349_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg465_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg2_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg7_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg372_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg563_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg226_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg101_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg516_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg182_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg516_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg562_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg265_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg562_out_to_MUX_Add3_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add3_3_impl_0_out);

   Delay1No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_3_impl_0_out,
                 Y => Delay1No58_out);

SharedReg589_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg589_out;
SharedReg424_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg424_out;
SharedReg151_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg151_out;
SharedReg122_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg122_out;
SharedReg698_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg698_out;
SharedReg181_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg181_out;
SharedReg347_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg347_out;
SharedReg653_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg653_out;
SharedReg267_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg267_out;
SharedReg656_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg656_out;
SharedReg18_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg18_out;
SharedReg23_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg23_out;
SharedReg425_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg425_out;
SharedReg511_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg511_out;
   MUX_Add3_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg589_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg424_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg18_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg23_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg425_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg511_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg151_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg122_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg698_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg181_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg347_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg653_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg267_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg656_out_to_MUX_Add3_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add3_3_impl_1_out);

   Delay1No59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_3_impl_1_out,
                 Y => Delay1No59_out);

Delay1No60_out_to_Add3_4_impl_parent_implementedSystem_port_0_cast <= Delay1No60_out;
Delay1No61_out_to_Add3_4_impl_parent_implementedSystem_port_1_cast <= Delay1No61_out;
   Add3_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add3_4_impl_out,
                 X => Delay1No60_out_to_Add3_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No61_out_to_Add3_4_impl_parent_implementedSystem_port_1_cast);

SharedReg302_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg302_out;
SharedReg568_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg568_out;
SharedReg356_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg356_out;
SharedReg469_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg469_out;
SharedReg234_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg234_out;
SharedReg104_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg104_out;
SharedReg523_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg523_out;
SharedReg190_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg190_out;
SharedReg523_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg523_out;
SharedReg567_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg567_out;
SharedReg274_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg274_out;
SharedReg567_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg567_out;
SharedReg2_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg2_out;
SharedReg7_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg7_out;
   MUX_Add3_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg302_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg568_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg274_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg567_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg2_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg7_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg356_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg469_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg234_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg104_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg523_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg190_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg523_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg567_out_to_MUX_Add3_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add3_4_impl_0_out);

   Delay1No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_4_impl_0_out,
                 Y => Delay1No60_out);

SharedReg448_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg448_out;
SharedReg518_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg518_out;
SharedReg594_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg594_out;
SharedReg392_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg392_out;
SharedReg156_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg156_out;
SharedReg127_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg127_out;
SharedReg703_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg703_out;
SharedReg189_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg189_out;
SharedReg354_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg354_out;
SharedReg658_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg658_out;
SharedReg276_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg276_out;
SharedReg661_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg661_out;
SharedReg18_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg18_out;
SharedReg23_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg23_out;
   MUX_Add3_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg448_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg518_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg276_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg661_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg18_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg23_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg594_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg392_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg156_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg127_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg703_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg189_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg354_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg658_out_to_MUX_Add3_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add3_4_impl_1_out);

   Delay1No61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add3_4_impl_1_out,
                 Y => Delay1No61_out);

Delay1No62_out_to_Add12_0_impl_parent_implementedSystem_port_0_cast <= Delay1No62_out;
Delay1No63_out_to_Add12_0_impl_parent_implementedSystem_port_1_cast <= Delay1No63_out;
   Add12_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_0_impl_out,
                 X => Delay1No62_out_to_Add12_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No63_out_to_Add12_0_impl_parent_implementedSystem_port_1_cast);

SharedReg198_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg198_out;
SharedReg3_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg3_out;
SharedReg8_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg8_out;
SharedReg377_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg377_out;
SharedReg239_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg239_out;
SharedReg134_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg134_out;
SharedReg283_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg283_out;
SharedReg303_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg303_out;
SharedReg132_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg132_out;
Delay10No60_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_10_cast <= Delay10No60_out;
SharedReg163_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg163_out;
SharedReg329_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg329_out;
SharedReg93_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg93_out;
SharedReg574_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg574_out;
   MUX_Add12_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg198_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg3_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg163_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg329_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg93_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg574_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg8_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg377_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg239_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg134_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg283_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg303_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg132_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay10No60_out_to_MUX_Add12_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add12_0_impl_0_out);

   Delay1No62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_0_impl_0_out,
                 Y => Delay1No62_out);

SharedReg243_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg243_out;
SharedReg19_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg24_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg24_out;
SharedReg394_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg394_out;
SharedReg157_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg157_out;
SharedReg237_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg237_out;
SharedReg450_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg450_out;
Delay4No75_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_8_cast <= Delay4No75_out;
SharedReg197_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg197_out;
Delay27No20_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_10_cast <= Delay27No20_out;
Delay28No_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_11_cast <= Delay28No_out;
SharedReg574_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg574_out;
SharedReg157_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg157_out;
SharedReg682_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg682_out;
   MUX_Add12_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg243_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay28No_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg574_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg157_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg682_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg24_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg394_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg157_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg237_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg450_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay4No75_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg197_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay27No20_out_to_MUX_Add12_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add12_0_impl_1_out);

   Delay1No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_0_impl_1_out,
                 Y => Delay1No63_out);

Delay1No64_out_to_Add12_1_impl_parent_implementedSystem_port_0_cast <= Delay1No64_out;
Delay1No65_out_to_Add12_1_impl_parent_implementedSystem_port_1_cast <= Delay1No65_out;
   Add12_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_1_impl_out,
                 X => Delay1No64_out_to_Add12_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No65_out_to_Add12_1_impl_parent_implementedSystem_port_1_cast);

SharedReg336_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg336_out;
SharedReg96_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg96_out;
SharedReg579_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg579_out;
SharedReg206_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg206_out;
SharedReg3_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg3_out;
SharedReg8_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg8_out;
SharedReg380_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg380_out;
SharedReg248_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg248_out;
SharedReg139_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg139_out;
SharedReg298_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg298_out;
SharedReg317_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg317_out;
SharedReg137_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg137_out;
Delay10No61_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_13_cast <= Delay10No61_out;
SharedReg171_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg171_out;
   MUX_Add12_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg336_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg96_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg317_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg137_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay10No61_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg171_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg579_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg206_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg3_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg8_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg380_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg248_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg139_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg298_out_to_MUX_Add12_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add12_1_impl_0_out);

   Delay1No64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_1_impl_0_out,
                 Y => Delay1No64_out);

SharedReg579_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg579_out;
SharedReg165_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg165_out;
SharedReg687_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg687_out;
SharedReg252_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg252_out;
SharedReg19_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg19_out;
SharedReg24_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg24_out;
SharedReg397_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg397_out;
SharedReg165_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg165_out;
SharedReg246_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg246_out;
SharedReg435_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg435_out;
Delay4No76_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_11_cast <= Delay4No76_out;
SharedReg205_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg205_out;
Delay27No21_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_13_cast <= Delay27No21_out;
Delay28No1_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_14_cast <= Delay28No1_out;
   MUX_Add12_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg579_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg165_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay4No76_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg205_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay27No21_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay28No1_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg687_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg252_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg19_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg24_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg397_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg165_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg246_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg435_out_to_MUX_Add12_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add12_1_impl_1_out);

   Delay1No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_1_impl_1_out,
                 Y => Delay1No65_out);

Delay1No66_out_to_Add12_2_impl_parent_implementedSystem_port_0_cast <= Delay1No66_out;
Delay1No67_out_to_Add12_2_impl_parent_implementedSystem_port_1_cast <= Delay1No67_out;
   Add12_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_2_impl_out,
                 X => Delay1No66_out_to_Add12_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No67_out_to_Add12_2_impl_parent_implementedSystem_port_1_cast);

SharedReg142_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg142_out;
Delay10No62_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_2_cast <= Delay10No62_out;
SharedReg179_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg179_out;
SharedReg343_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg343_out;
SharedReg99_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg99_out;
SharedReg584_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg584_out;
SharedReg214_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg214_out;
SharedReg3_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg3_out;
SharedReg8_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg8_out;
SharedReg401_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg401_out;
SharedReg257_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg257_out;
SharedReg144_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg144_out;
SharedReg308_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg308_out;
SharedReg367_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg367_out;
   MUX_Add12_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg142_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay10No62_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg257_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg144_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg308_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg367_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg179_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg343_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg99_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg584_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg214_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg3_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg8_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg401_out_to_MUX_Add12_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add12_2_impl_0_out);

   Delay1No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_2_impl_0_out,
                 Y => Delay1No66_out);

SharedReg213_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg213_out;
Delay27No22_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_2_cast <= Delay27No22_out;
Delay28No2_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_3_cast <= Delay28No2_out;
SharedReg584_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg584_out;
SharedReg173_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg173_out;
SharedReg692_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg692_out;
SharedReg261_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg261_out;
SharedReg19_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg19_out;
SharedReg24_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg24_out;
SharedReg419_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg419_out;
SharedReg173_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg173_out;
SharedReg255_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg255_out;
SharedReg457_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg457_out;
SharedReg385_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg385_out;
   MUX_Add12_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg213_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay27No22_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg173_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg255_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg457_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg385_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => Delay28No2_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg584_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg173_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg692_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg261_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg19_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg24_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg419_out_to_MUX_Add12_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add12_2_impl_1_out);

   Delay1No67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_2_impl_1_out,
                 Y => Delay1No67_out);

Delay1No68_out_to_Add12_3_impl_parent_implementedSystem_port_0_cast <= Delay1No68_out;
Delay1No69_out_to_Add12_3_impl_parent_implementedSystem_port_1_cast <= Delay1No69_out;
   Add12_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_3_impl_out,
                 X => Delay1No68_out_to_Add12_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No69_out_to_Add12_3_impl_parent_implementedSystem_port_1_cast);

SharedReg149_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg149_out;
SharedReg313_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg313_out;
SharedReg312_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg312_out;
SharedReg147_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg147_out;
Delay10No63_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_5_cast <= Delay10No63_out;
SharedReg187_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg187_out;
SharedReg350_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg350_out;
SharedReg102_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg102_out;
SharedReg589_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg589_out;
SharedReg222_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg222_out;
SharedReg3_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg3_out;
SharedReg8_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg8_out;
SharedReg404_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg404_out;
SharedReg266_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg266_out;
   MUX_Add12_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg149_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg313_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg3_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg8_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg404_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg266_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg312_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg147_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay10No63_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg187_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg350_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg102_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg589_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg222_out_to_MUX_Add12_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add12_3_impl_0_out);

   Delay1No68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_3_impl_0_out,
                 Y => Delay1No68_out);

SharedReg264_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg264_out;
SharedReg443_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg443_out;
SharedReg389_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg389_out;
SharedReg221_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg221_out;
Delay27No23_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_5_cast <= Delay27No23_out;
Delay28No3_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_6_cast <= Delay28No3_out;
SharedReg589_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg589_out;
SharedReg181_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg181_out;
SharedReg697_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg697_out;
SharedReg270_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg270_out;
SharedReg19_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg19_out;
SharedReg24_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg24_out;
SharedReg423_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg423_out;
SharedReg181_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg181_out;
   MUX_Add12_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg264_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg443_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg19_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg24_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg423_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg181_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg389_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg221_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay27No23_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay28No3_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg589_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg181_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg697_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg270_out_to_MUX_Add12_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add12_3_impl_1_out);

   Delay1No69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_3_impl_1_out,
                 Y => Delay1No69_out);

Delay1No70_out_to_Add12_4_impl_parent_implementedSystem_port_0_cast <= Delay1No70_out;
Delay1No71_out_to_Add12_4_impl_parent_implementedSystem_port_1_cast <= Delay1No71_out;
   Add12_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add12_4_impl_out,
                 X => Delay1No70_out_to_Add12_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No71_out_to_Add12_4_impl_parent_implementedSystem_port_1_cast);

SharedReg408_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg408_out;
SharedReg275_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg275_out;
SharedReg154_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg154_out;
SharedReg301_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg301_out;
SharedReg300_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg300_out;
SharedReg152_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg152_out;
Delay10No64_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_7_cast <= Delay10No64_out;
SharedReg195_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg195_out;
SharedReg357_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg357_out;
SharedReg105_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg105_out;
SharedReg594_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg594_out;
SharedReg230_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg230_out;
SharedReg3_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg3_out;
SharedReg8_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg8_out;
   MUX_Add12_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg408_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg275_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg594_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg230_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg3_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg8_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg154_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg301_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg300_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg152_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay10No64_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg195_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg357_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg105_out_to_MUX_Add12_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add12_4_impl_0_out);

   Delay1No70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_4_impl_0_out,
                 Y => Delay1No70_out);

SharedReg427_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg427_out;
SharedReg189_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg189_out;
SharedReg273_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg273_out;
SharedReg466_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg466_out;
SharedReg324_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg324_out;
SharedReg229_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg229_out;
Delay27No24_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_7_cast <= Delay27No24_out;
Delay28No4_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_8_cast <= Delay28No4_out;
SharedReg594_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg594_out;
SharedReg189_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg189_out;
SharedReg702_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg702_out;
SharedReg279_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg279_out;
SharedReg19_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg19_out;
SharedReg24_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg24_out;
   MUX_Add12_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg427_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg189_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg702_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg279_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg19_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg24_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg273_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg466_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg324_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg229_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay27No24_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay28No4_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg594_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg189_out_to_MUX_Add12_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add12_4_impl_1_out);

   Delay1No71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add12_4_impl_1_out,
                 Y => Delay1No71_out);

Delay1No72_out_to_Add9_0_impl_parent_implementedSystem_port_0_cast <= Delay1No72_out;
Delay1No73_out_to_Add9_0_impl_parent_implementedSystem_port_1_cast <= Delay1No73_out;
   Add9_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add9_0_impl_out,
                 X => Delay1No72_out_to_Add9_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No73_out_to_Add9_0_impl_parent_implementedSystem_port_1_cast);

SharedReg238_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg238_out;
SharedReg4_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg4_out;
SharedReg9_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg9_out;
SharedReg395_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg395_out;
SharedReg326_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg326_out;
SharedReg453_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg453_out;
SharedReg411_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg411_out;
SharedReg305_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg305_out;
SharedReg362_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg362_out;
SharedReg245_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg245_out;
SharedReg495_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg495_out;
SharedReg376_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg376_out;
SharedReg546_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg546_out;
SharedReg361_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg361_out;
   MUX_Add9_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg238_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg4_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg495_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg376_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg546_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg361_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg9_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg395_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg326_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg453_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg411_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg305_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg362_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg245_out_to_MUX_Add9_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add9_0_impl_0_out);

   Delay1No72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_0_impl_0_out,
                 Y => Delay1No72_out);

SharedReg242_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg242_out;
SharedReg20_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg25_out;
SharedReg412_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg412_out;
SharedReg547_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg547_out;
SharedReg431_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg431_out;
SharedReg431_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg431_out;
SharedReg528_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg528_out;
SharedReg282_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg282_out;
Delay27No15_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_10_cast <= Delay27No15_out;
SharedReg743_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg743_out;
SharedReg393_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg393_out;
SharedReg493_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg493_out;
SharedReg376_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg376_out;
   MUX_Add9_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg242_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg743_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg393_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg493_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg376_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg25_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg412_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg547_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg431_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg431_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg528_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg282_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay27No15_out_to_MUX_Add9_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add9_0_impl_1_out);

   Delay1No73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_0_impl_1_out,
                 Y => Delay1No73_out);

Delay1No74_out_to_Add9_1_impl_parent_implementedSystem_port_0_cast <= Delay1No74_out;
Delay1No75_out_to_Add9_1_impl_parent_implementedSystem_port_1_cast <= Delay1No75_out;
   Add9_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add9_1_impl_out,
                 X => Delay1No74_out_to_Add9_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No75_out_to_Add9_1_impl_parent_implementedSystem_port_1_cast);

SharedReg379_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg379_out;
SharedReg551_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg551_out;
SharedReg317_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg317_out;
SharedReg247_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg247_out;
SharedReg4_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg4_out;
SharedReg9_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg9_out;
SharedReg398_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg398_out;
SharedReg333_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg333_out;
SharedReg456_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg456_out;
SharedReg415_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg415_out;
SharedReg319_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg319_out;
SharedReg365_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg365_out;
SharedReg254_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg254_out;
SharedReg502_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg502_out;
   MUX_Add9_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg379_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg551_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg319_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg365_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg254_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg502_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg317_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg247_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg4_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg9_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg398_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg333_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg456_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg415_out_to_MUX_Add9_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add9_1_impl_0_out);

   Delay1No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_1_impl_0_out,
                 Y => Delay1No74_out);

SharedReg396_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg396_out;
SharedReg500_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg500_out;
SharedReg364_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg364_out;
SharedReg251_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg251_out;
SharedReg20_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg25_out;
SharedReg416_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg416_out;
SharedReg552_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg552_out;
SharedReg436_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg436_out;
SharedReg436_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg436_out;
SharedReg533_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg533_out;
SharedReg297_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg297_out;
Delay27No16_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_13_cast <= Delay27No16_out;
SharedReg751_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg751_out;
   MUX_Add9_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg396_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg500_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg533_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg297_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay27No16_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg751_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg364_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg251_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg20_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg25_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg416_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg552_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg436_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg436_out_to_MUX_Add9_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add9_1_impl_1_out);

   Delay1No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_1_impl_1_out,
                 Y => Delay1No75_out);

Delay1No76_out_to_Add9_2_impl_parent_implementedSystem_port_0_cast <= Delay1No76_out;
Delay1No77_out_to_Add9_2_impl_parent_implementedSystem_port_1_cast <= Delay1No77_out;
   Add9_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add9_2_impl_out,
                 X => Delay1No76_out_to_Add9_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No77_out_to_Add9_2_impl_parent_implementedSystem_port_1_cast);

SharedReg383_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg383_out;
SharedReg263_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg263_out;
SharedReg509_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg509_out;
SharedReg382_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg382_out;
SharedReg556_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg556_out;
SharedReg367_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg367_out;
SharedReg256_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg256_out;
SharedReg4_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg4_out;
SharedReg9_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg9_out;
SharedReg420_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg420_out;
SharedReg340_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg340_out;
SharedReg481_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg481_out;
SharedReg440_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg440_out;
SharedReg369_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg369_out;
   MUX_Add9_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg383_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg263_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg340_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg481_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg440_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg369_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg509_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg382_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg556_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg367_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg256_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg4_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg9_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg420_out_to_MUX_Add9_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add9_2_impl_0_out);

   Delay1No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_2_impl_0_out,
                 Y => Delay1No76_out);

SharedReg307_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg307_out;
Delay27No17_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_2_cast <= Delay27No17_out;
SharedReg759_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg759_out;
SharedReg400_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg400_out;
SharedReg507_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg507_out;
SharedReg382_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg382_out;
SharedReg260_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg260_out;
SharedReg20_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg25_out;
SharedReg441_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg441_out;
SharedReg557_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg557_out;
SharedReg458_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg458_out;
SharedReg458_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg458_out;
SharedReg603_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg603_out;
   MUX_Add9_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg307_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay27No17_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg557_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg458_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg458_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg603_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg759_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg400_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg507_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg382_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg260_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg20_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg25_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg441_out_to_MUX_Add9_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add9_2_impl_1_out);

   Delay1No77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_2_impl_1_out,
                 Y => Delay1No77_out);

Delay1No78_out_to_Add9_3_impl_parent_implementedSystem_port_0_cast <= Delay1No78_out;
Delay1No79_out_to_Add9_3_impl_parent_implementedSystem_port_1_cast <= Delay1No79_out;
   Add9_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add9_3_impl_out,
                 X => Delay1No78_out_to_Add9_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No79_out_to_Add9_3_impl_parent_implementedSystem_port_1_cast);

SharedReg485_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg485_out;
SharedReg444_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg444_out;
SharedReg372_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg372_out;
SharedReg371_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg371_out;
SharedReg272_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg272_out;
SharedReg516_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg516_out;
SharedReg386_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg386_out;
SharedReg561_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg561_out;
SharedReg370_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg370_out;
SharedReg265_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg265_out;
SharedReg4_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg4_out;
SharedReg9_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg9_out;
SharedReg424_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg424_out;
SharedReg347_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg347_out;
   MUX_Add9_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg485_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg444_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg4_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg9_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg424_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg347_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg372_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg371_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg272_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg516_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg386_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg561_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg370_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg265_out_to_MUX_Add9_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add9_3_impl_0_out);

   Delay1No78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_3_impl_0_out,
                 Y => Delay1No78_out);

SharedReg462_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg462_out;
SharedReg462_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg462_out;
SharedReg609_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg609_out;
SharedReg292_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg292_out;
Delay27No18_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_5_cast <= Delay27No18_out;
SharedReg767_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg767_out;
SharedReg403_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg403_out;
SharedReg514_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg514_out;
SharedReg386_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg386_out;
SharedReg269_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg269_out;
SharedReg20_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg25_out;
SharedReg445_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg445_out;
SharedReg562_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg562_out;
   MUX_Add9_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg462_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg462_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg20_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg25_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg445_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg609_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg292_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay27No18_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg767_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg403_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg514_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg386_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg269_out_to_MUX_Add9_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add9_3_impl_1_out);

   Delay1No79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_3_impl_1_out,
                 Y => Delay1No79_out);

Delay1No80_out_to_Add9_4_impl_parent_implementedSystem_port_0_cast <= Delay1No80_out;
Delay1No81_out_to_Add9_4_impl_parent_implementedSystem_port_1_cast <= Delay1No81_out;
   Add9_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add9_4_impl_out,
                 X => Delay1No80_out_to_Add9_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No81_out_to_Add9_4_impl_parent_implementedSystem_port_1_cast);

SharedReg392_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg392_out;
SharedReg354_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg354_out;
SharedReg449_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg449_out;
SharedReg427_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg427_out;
SharedReg323_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg323_out;
SharedReg322_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg322_out;
SharedReg281_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg281_out;
SharedReg523_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg523_out;
SharedReg390_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg390_out;
SharedReg566_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg566_out;
SharedReg373_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg373_out;
SharedReg274_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg274_out;
SharedReg4_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg4_out;
SharedReg9_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg9_out;
   MUX_Add9_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg392_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg354_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg373_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg274_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg4_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg9_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg449_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg427_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg323_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg322_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg281_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg523_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg390_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg566_out_to_MUX_Add9_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add9_4_impl_0_out);

   Delay1No80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_4_impl_0_out,
                 Y => Delay1No80_out);

SharedReg409_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg409_out;
SharedReg567_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg567_out;
SharedReg427_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg427_out;
SharedReg447_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg447_out;
SharedReg614_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg614_out;
SharedReg300_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg300_out;
Delay27No19_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_7_cast <= Delay27No19_out;
SharedReg775_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg775_out;
SharedReg407_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg407_out;
SharedReg521_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg521_out;
SharedReg390_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg390_out;
SharedReg278_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg278_out;
SharedReg20_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg20_out;
SharedReg25_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg25_out;
   MUX_Add9_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg409_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg567_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg390_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg278_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg20_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg25_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg427_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg447_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg614_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg300_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay27No19_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg775_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg407_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg521_out_to_MUX_Add9_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add9_4_impl_1_out);

   Delay1No81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add9_4_impl_1_out,
                 Y => Delay1No81_out);

Delay1No82_out_to_Add18_0_impl_parent_implementedSystem_port_0_cast <= Delay1No82_out;
Delay1No83_out_to_Add18_0_impl_parent_implementedSystem_port_1_cast <= Delay1No83_out;
   Add18_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add18_0_impl_out,
                 X => Delay1No82_out_to_Add18_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No83_out_to_Add18_0_impl_parent_implementedSystem_port_1_cast);

SharedReg361_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg361_out;
SharedReg5_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg10_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg10_out;
SharedReg472_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg472_out;
SharedReg132_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg132_out;
SharedReg527_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg527_out;
SharedReg526_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg526_out;
SharedReg526_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg526_out;
SharedReg376_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg376_out;
Delay15No10_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_10_cast <= Delay15No10_out;
SharedReg245_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg245_out;
SharedReg283_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg283_out;
SharedReg283_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg283_out;
SharedReg393_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg393_out;
   MUX_Add18_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg361_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg245_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg283_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg283_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg393_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg10_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg472_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg132_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg527_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg526_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg526_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg376_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay15No10_out_to_MUX_Add18_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add18_0_impl_0_out);

   Delay1No82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_0_impl_0_out,
                 Y => Delay1No82_out);

SharedReg376_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg376_out;
SharedReg21_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg21_out;
SharedReg26_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg26_out;
SharedReg473_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg473_out;
SharedReg238_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg238_out;
SharedReg526_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg526_out;
SharedReg617_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg617_out;
SharedReg617_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg617_out;
SharedReg393_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg393_out;
SharedReg361_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg361_out;
SharedReg204_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg204_out;
SharedReg450_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg450_out;
SharedReg303_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg303_out;
SharedReg451_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg451_out;
   MUX_Add18_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg376_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg21_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg204_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg450_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg303_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg451_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg26_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg473_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg238_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg526_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg617_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg617_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg393_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg361_out_to_MUX_Add18_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add18_0_impl_1_out);

   Delay1No83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_0_impl_1_out,
                 Y => Delay1No83_out);

Delay1No84_out_to_Add18_1_impl_parent_implementedSystem_port_0_cast <= Delay1No84_out;
Delay1No85_out_to_Add18_1_impl_parent_implementedSystem_port_1_cast <= Delay1No85_out;
   Add18_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add18_1_impl_out,
                 X => Delay1No84_out_to_Add18_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No85_out_to_Add18_1_impl_parent_implementedSystem_port_1_cast);

SharedReg298_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg298_out;
SharedReg298_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg298_out;
SharedReg379_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg379_out;
SharedReg317_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg317_out;
SharedReg5_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg5_out;
SharedReg10_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg10_out;
SharedReg477_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg477_out;
SharedReg137_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg137_out;
SharedReg532_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg532_out;
SharedReg530_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg530_out;
SharedReg476_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg476_out;
SharedReg379_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg379_out;
Delay15No11_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_13_cast <= Delay15No11_out;
SharedReg254_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg254_out;
   MUX_Add18_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg298_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg298_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg476_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg379_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay15No11_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg254_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg379_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg317_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg5_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg10_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg477_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg137_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg532_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg530_out_to_MUX_Add18_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add18_1_impl_0_out);

   Delay1No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_1_impl_0_out,
                 Y => Delay1No84_out);

SharedReg454_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg454_out;
SharedReg297_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg297_out;
SharedReg436_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg436_out;
SharedReg364_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg364_out;
SharedReg21_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg21_out;
SharedReg26_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg26_out;
SharedReg455_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg455_out;
SharedReg247_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg247_out;
SharedReg530_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg530_out;
SharedReg622_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg622_out;
SharedReg530_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg530_out;
SharedReg396_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg396_out;
SharedReg364_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg364_out;
SharedReg212_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg212_out;
   MUX_Add18_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg454_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg297_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg530_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg396_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg364_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg212_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg436_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg364_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg21_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg26_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg455_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg247_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg530_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg622_out_to_MUX_Add18_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add18_1_impl_1_out);

   Delay1No85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_1_impl_1_out,
                 Y => Delay1No85_out);

Delay1No86_out_to_Add18_2_impl_parent_implementedSystem_port_0_cast <= Delay1No86_out;
Delay1No87_out_to_Add18_2_impl_parent_implementedSystem_port_1_cast <= Delay1No87_out;
   Add18_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add18_2_impl_out,
                 X => Delay1No86_out_to_Add18_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No87_out_to_Add18_2_impl_parent_implementedSystem_port_1_cast);

SharedReg400_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg400_out;
Delay15No12_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_2_cast <= Delay15No12_out;
SharedReg263_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg263_out;
SharedReg290_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg290_out;
SharedReg290_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg290_out;
SharedReg400_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg400_out;
SharedReg367_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg367_out;
SharedReg5_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg5_out;
SharedReg10_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg10_out;
SharedReg536_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg536_out;
SharedReg142_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg142_out;
SharedReg602_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg602_out;
SharedReg600_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg600_out;
SharedReg535_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg535_out;
   MUX_Add18_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg400_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay15No12_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg142_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg602_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg600_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg535_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg263_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg290_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg290_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg400_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg367_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg5_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg10_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg536_out_to_MUX_Add18_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add18_2_impl_0_out);

   Delay1No86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_2_impl_0_out,
                 Y => Delay1No86_out);

SharedReg418_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg418_out;
SharedReg367_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg367_out;
SharedReg220_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg220_out;
SharedReg457_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg457_out;
SharedReg307_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg307_out;
SharedReg458_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg458_out;
SharedReg382_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg382_out;
SharedReg21_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg21_out;
SharedReg26_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg26_out;
SharedReg480_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg480_out;
SharedReg256_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg256_out;
SharedReg600_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg600_out;
SharedReg627_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg627_out;
SharedReg600_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg600_out;
   MUX_Add18_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg418_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg367_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg256_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg600_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg627_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg600_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg220_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg457_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg307_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg458_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg382_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg21_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg26_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg480_out_to_MUX_Add18_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add18_2_impl_1_out);

   Delay1No87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_2_impl_1_out,
                 Y => Delay1No87_out);

Delay1No88_out_to_Add18_3_impl_parent_implementedSystem_port_0_cast <= Delay1No88_out;
Delay1No89_out_to_Add18_3_impl_parent_implementedSystem_port_1_cast <= Delay1No89_out;
   Add18_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add18_3_impl_out,
                 X => Delay1No88_out_to_Add18_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No89_out_to_Add18_3_impl_parent_implementedSystem_port_1_cast);

SharedReg608_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg608_out;
SharedReg606_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg606_out;
SharedReg483_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg483_out;
SharedReg386_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg386_out;
Delay15No13_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_5_cast <= Delay15No13_out;
SharedReg272_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg272_out;
SharedReg293_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg293_out;
SharedReg293_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg293_out;
SharedReg403_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg403_out;
SharedReg312_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg312_out;
SharedReg5_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg5_out;
SharedReg10_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg10_out;
SharedReg540_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg540_out;
SharedReg147_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg147_out;
   MUX_Add18_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg608_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg606_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg5_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg10_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg540_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg147_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg483_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg386_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay15No13_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg272_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg293_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg293_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg403_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg312_out_to_MUX_Add18_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add18_3_impl_0_out);

   Delay1No88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_3_impl_0_out,
                 Y => Delay1No88_out);

SharedReg606_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg606_out;
SharedReg630_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg630_out;
SharedReg539_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg539_out;
SharedReg403_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg403_out;
SharedReg370_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg370_out;
SharedReg228_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg228_out;
SharedReg461_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg461_out;
SharedReg312_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg312_out;
SharedReg462_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg462_out;
SharedReg370_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg370_out;
SharedReg21_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg21_out;
SharedReg26_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg26_out;
SharedReg464_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg464_out;
SharedReg265_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg265_out;
   MUX_Add18_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg606_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg630_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg21_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg26_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg464_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg265_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg539_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg403_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg370_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg228_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg461_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg312_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg462_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg370_out_to_MUX_Add18_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add18_3_impl_1_out);

   Delay1No89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_3_impl_1_out,
                 Y => Delay1No89_out);

Delay1No90_out_to_Add18_4_impl_parent_implementedSystem_port_0_cast <= Delay1No90_out;
Delay1No91_out_to_Add18_4_impl_parent_implementedSystem_port_1_cast <= Delay1No91_out;
   Add18_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add18_4_impl_out,
                 X => Delay1No90_out_to_Add18_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No91_out_to_Add18_4_impl_parent_implementedSystem_port_1_cast);

SharedReg468_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg468_out;
SharedReg152_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg152_out;
SharedReg489_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg489_out;
SharedReg543_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg543_out;
SharedReg543_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg543_out;
SharedReg390_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg390_out;
Delay15No14_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_7_cast <= Delay15No14_out;
SharedReg281_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg281_out;
SharedReg301_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg301_out;
SharedReg301_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg301_out;
SharedReg407_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg407_out;
SharedReg373_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg373_out;
SharedReg5_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg5_out;
SharedReg10_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg10_out;
   MUX_Add18_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg468_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg152_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg407_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg373_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg5_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg10_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg489_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg543_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg543_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg390_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay15No14_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg281_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg301_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg301_out_to_MUX_Add18_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add18_4_impl_0_out);

   Delay1No90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_4_impl_0_out,
                 Y => Delay1No90_out);

SharedReg488_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg488_out;
SharedReg274_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg274_out;
SharedReg487_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg487_out;
SharedReg612_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg612_out;
SharedReg612_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg612_out;
SharedReg407_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg407_out;
SharedReg373_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg373_out;
SharedReg236_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg236_out;
SharedReg466_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg466_out;
SharedReg300_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg300_out;
SharedReg447_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg447_out;
SharedReg390_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg390_out;
SharedReg21_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg21_out;
SharedReg26_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg26_out;
   MUX_Add18_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg488_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg274_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg447_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg390_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg21_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg26_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg487_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg612_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg612_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg407_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg373_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg236_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg466_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg300_out_to_MUX_Add18_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add18_4_impl_1_out);

   Delay1No91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add18_4_impl_1_out,
                 Y => Delay1No91_out);

Delay1No92_out_to_Add128_0_impl_parent_implementedSystem_port_0_cast <= Delay1No92_out;
Delay1No93_out_to_Add128_0_impl_parent_implementedSystem_port_1_cast <= Delay1No93_out;
   Add128_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add128_0_impl_out,
                 X => Delay1No92_out_to_Add128_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No93_out_to_Add128_0_impl_parent_implementedSystem_port_1_cast);

SharedReg618_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg618_out;
SharedReg13_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg13_out;
SharedReg11_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg11_out;
SharedReg617_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg617_out;
SharedReg285_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg285_out;
SharedReg617_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg617_out;
SharedReg671_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg671_out;
SharedReg430_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg430_out;
SharedReg377_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg377_out;
SharedReg471_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg471_out;
SharedReg410_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg410_out;
SharedReg632_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg632_out;
SharedReg376_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg376_out;
SharedReg450_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg450_out;
   MUX_Add128_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg618_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg410_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg632_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg376_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg450_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg11_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg617_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg285_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg617_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg671_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg430_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg377_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg471_out_to_MUX_Add128_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add128_0_impl_0_out);

   Delay1No92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_0_impl_0_out,
                 Y => Delay1No92_out);

SharedReg632_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg632_out;
SharedReg29_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg29_out;
SharedReg27_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg27_out;
SharedReg672_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg672_out;
SharedReg305_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg305_out;
SharedReg305_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg305_out;
SharedReg286_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg286_out;
SharedReg450_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg450_out;
SharedReg450_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg450_out;
Delay15No25_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_10_cast <= Delay15No25_out;
SharedReg430_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg430_out;
SharedReg617_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg617_out;
SharedReg393_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg393_out;
SharedReg470_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg470_out;
   MUX_Add128_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg632_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg29_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg430_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg617_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg393_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg470_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg27_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg672_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg305_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg305_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg286_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg450_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg450_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay15No25_out_to_MUX_Add128_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add128_0_impl_1_out);

   Delay1No93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_0_impl_1_out,
                 Y => Delay1No93_out);

Delay1No94_out_to_Add128_1_impl_parent_implementedSystem_port_0_cast <= Delay1No94_out;
Delay1No95_out_to_Add128_1_impl_parent_implementedSystem_port_1_cast <= Delay1No95_out;
   Add128_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add128_1_impl_out,
                 X => Delay1No94_out_to_Add128_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No95_out_to_Add128_1_impl_parent_implementedSystem_port_1_cast);

SharedReg662_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg662_out;
SharedReg364_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg364_out;
SharedReg435_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg435_out;
SharedReg531_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg531_out;
SharedReg13_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg13_out;
SharedReg11_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg11_out;
SharedReg622_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg622_out;
Delay4No71_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_8_cast <= Delay4No71_out;
SharedReg622_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg622_out;
SharedReg674_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg674_out;
SharedReg435_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg435_out;
SharedReg380_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg380_out;
SharedReg476_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg476_out;
SharedReg414_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg414_out;
   MUX_Add128_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg662_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg364_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg435_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg380_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg476_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg414_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg435_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg531_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg13_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg11_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg622_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay4No71_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg622_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg674_out_to_MUX_Add128_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add128_1_impl_0_out);

   Delay1No94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_1_impl_0_out,
                 Y => Delay1No94_out);

SharedReg622_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg622_out;
SharedReg379_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg379_out;
SharedReg454_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg454_out;
SharedReg621_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg621_out;
SharedReg29_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg29_out;
SharedReg27_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg27_out;
SharedReg675_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg675_out;
SharedReg319_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg319_out;
SharedReg319_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg319_out;
SharedReg673_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg673_out;
SharedReg454_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg454_out;
SharedReg454_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg454_out;
Delay15No26_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_13_cast <= Delay15No26_out;
SharedReg435_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg435_out;
   MUX_Add128_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg622_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg379_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg454_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg454_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay15No26_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg435_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg454_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg621_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg29_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg27_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg675_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg319_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg319_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg673_out_to_MUX_Add128_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add128_1_impl_1_out);

   Delay1No95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_1_impl_1_out,
                 Y => Delay1No95_out);

Delay1No96_out_to_Add128_2_impl_parent_implementedSystem_port_0_cast <= Delay1No96_out;
Delay1No97_out_to_Add128_2_impl_parent_implementedSystem_port_1_cast <= Delay1No97_out;
   Add128_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add128_2_impl_out,
                 X => Delay1No96_out_to_Add128_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No97_out_to_Add128_2_impl_parent_implementedSystem_port_1_cast);

SharedReg401_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg401_out;
SharedReg535_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg535_out;
SharedReg418_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg418_out;
SharedReg626_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg626_out;
SharedReg382_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg382_out;
SharedReg457_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg457_out;
SharedReg601_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg601_out;
SharedReg13_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg13_out;
SharedReg11_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg11_out;
SharedReg627_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg627_out;
SharedReg310_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg310_out;
SharedReg627_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg627_out;
SharedReg572_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg572_out;
SharedReg457_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg457_out;
   MUX_Add128_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg401_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg535_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg310_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg627_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg572_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg457_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg418_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg626_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg382_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg457_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg601_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg13_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg11_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg627_out_to_MUX_Add128_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add128_2_impl_0_out);

   Delay1No96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_2_impl_0_out,
                 Y => Delay1No96_out);

SharedReg479_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg479_out;
Delay15No27_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_2_cast <= Delay15No27_out;
SharedReg439_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg439_out;
SharedReg600_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg600_out;
SharedReg400_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg400_out;
SharedReg479_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg479_out;
SharedReg626_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg626_out;
SharedReg29_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg29_out;
SharedReg27_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg27_out;
SharedReg573_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg573_out;
SharedReg369_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg369_out;
SharedReg309_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg309_out;
SharedReg571_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg571_out;
SharedReg479_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg479_out;
   MUX_Add128_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg479_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay15No27_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg369_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg309_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg571_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg479_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg439_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg600_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg400_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg479_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg626_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg29_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg27_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg573_out_to_MUX_Add128_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add128_2_impl_1_out);

   Delay1No97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_2_impl_1_out,
                 Y => Delay1No97_out);

Delay1No98_out_to_Add128_3_impl_parent_implementedSystem_port_0_cast <= Delay1No98_out;
Delay1No99_out_to_Add128_3_impl_parent_implementedSystem_port_1_cast <= Delay1No99_out;
   Add128_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add128_3_impl_out,
                 X => Delay1No98_out_to_Add128_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No99_out_to_Add128_3_impl_parent_implementedSystem_port_1_cast);

SharedReg630_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg630_out;
SharedReg295_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg295_out;
SharedReg443_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg443_out;
SharedReg387_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg387_out;
SharedReg483_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg483_out;
SharedReg422_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg422_out;
SharedReg629_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg629_out;
SharedReg386_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg386_out;
SharedReg461_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg461_out;
SharedReg607_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg607_out;
SharedReg13_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg13_out;
SharedReg11_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg11_out;
SharedReg630_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg630_out;
SharedReg315_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg315_out;
   MUX_Add128_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg630_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg295_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg13_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg11_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg630_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg315_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg443_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg387_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg483_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg422_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg629_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg386_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg461_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg607_out_to_MUX_Add128_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add128_3_impl_0_out);

   Delay1No98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_3_impl_0_out,
                 Y => Delay1No98_out);

SharedReg314_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg314_out;
SharedReg667_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg667_out;
SharedReg461_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg461_out;
SharedReg461_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg461_out;
Delay15No28_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_5_cast <= Delay15No28_out;
SharedReg443_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg443_out;
SharedReg606_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg606_out;
SharedReg403_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg403_out;
SharedReg482_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg482_out;
SharedReg605_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg605_out;
SharedReg29_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg29_out;
SharedReg27_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg27_out;
SharedReg296_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg296_out;
SharedReg372_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg372_out;
   MUX_Add128_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg314_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg667_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg29_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg27_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg296_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg372_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg461_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg461_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay15No28_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg443_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg606_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg403_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg482_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg605_out_to_MUX_Add128_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add128_3_impl_1_out);

   Delay1No99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_3_impl_1_out,
                 Y => Delay1No99_out);

Delay1No100_out_to_Add128_4_impl_parent_implementedSystem_port_0_cast <= Delay1No100_out;
Delay1No101_out_to_Add128_4_impl_parent_implementedSystem_port_1_cast <= Delay1No101_out;
   Add128_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add128_4_impl_out,
                 X => Delay1No100_out_to_Add128_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No101_out_to_Add128_4_impl_parent_implementedSystem_port_1_cast);

SharedReg636_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg636_out;
Delay4No74_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_2_cast <= Delay4No74_out;
SharedReg543_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg543_out;
SharedReg677_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg677_out;
SharedReg426_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg426_out;
SharedReg374_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg374_out;
SharedReg487_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg487_out;
SharedReg426_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg426_out;
SharedReg635_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg635_out;
SharedReg373_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg373_out;
SharedReg466_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg466_out;
SharedReg544_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg544_out;
SharedReg13_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg13_out;
SharedReg11_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg11_out;
   MUX_Add128_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg636_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay4No74_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg466_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg544_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg13_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg11_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg543_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg677_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg426_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg374_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg487_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg426_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg635_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg373_out_to_MUX_Add128_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add128_4_impl_0_out);

   Delay1No100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_4_impl_0_out,
                 Y => Delay1No100_out);

Delay3No214_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_1_cast <= Delay3No214_out;
SharedReg375_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg375_out;
SharedReg375_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg375_out;
SharedReg734_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg734_out;
SharedReg446_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg446_out;
SharedReg466_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg466_out;
Delay15No29_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_7_cast <= Delay15No29_out;
SharedReg446_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg446_out;
SharedReg612_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg612_out;
SharedReg390_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg390_out;
SharedReg486_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg486_out;
SharedReg635_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg635_out;
SharedReg29_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg29_out;
SharedReg27_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg27_out;
   MUX_Add128_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay3No214_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg375_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg486_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg635_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg29_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg27_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg375_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg734_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg446_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg466_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay15No29_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg446_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg612_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg390_out_to_MUX_Add128_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add128_4_impl_1_out);

   Delay1No101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add128_4_impl_1_out,
                 Y => Delay1No101_out);

Delay1No102_out_to_Add40_0_impl_parent_implementedSystem_port_0_cast <= Delay1No102_out;
Delay1No103_out_to_Add40_0_impl_parent_implementedSystem_port_1_cast <= Delay1No103_out;
   Add40_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add40_0_impl_out,
                 X => Delay1No102_out_to_Add40_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No103_out_to_Add40_0_impl_parent_implementedSystem_port_1_cast);

SharedReg617_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg617_out;
SharedReg15_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg15_out;
SharedReg14_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg14_out;
SharedReg430_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg430_out;
SharedReg617_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg617_out;
SharedReg633_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg633_out;
Delay11No30_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_7_cast <= Delay11No30_out;
SharedReg525_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg525_out;
SharedReg671_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg671_out;
SharedReg617_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg617_out;
Delay16No_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_11_cast <= Delay16No_out;
SharedReg287_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg287_out;
SharedReg363_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg363_out;
SharedReg286_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg286_out;
   MUX_Add40_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg617_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay16No_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg287_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg363_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg286_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg14_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg430_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg617_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg633_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay11No30_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg525_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg671_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg617_out_to_MUX_Add40_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add40_0_impl_0_out);

   Delay1No102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_0_impl_0_out,
                 Y => Delay1No102_out);

SharedReg286_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg286_out;
SharedReg31_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg31_out;
SharedReg30_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg30_out;
SharedReg450_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg450_out;
SharedReg633_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg633_out;
SharedReg395_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg395_out;
SharedReg288_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg288_out;
SharedReg616_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg616_out;
SharedReg286_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg286_out;
Delay15No35_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_10_cast <= Delay15No35_out;
SharedReg633_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg633_out;
SharedReg670_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg670_out;
SharedReg525_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg525_out;
SharedReg671_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg671_out;
   MUX_Add40_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg286_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg31_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg633_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg670_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg525_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg671_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg30_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg450_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg633_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg395_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg288_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg616_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg286_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay15No35_out_to_MUX_Add40_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add40_0_impl_1_out);

   Delay1No103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_0_impl_1_out,
                 Y => Delay1No103_out);

Delay1No104_out_to_Add40_1_impl_parent_implementedSystem_port_0_cast <= Delay1No104_out;
Delay1No105_out_to_Add40_1_impl_parent_implementedSystem_port_1_cast <= Delay1No105_out;
   Add40_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add40_1_impl_out,
                 X => Delay1No104_out_to_Add40_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No105_out_to_Add40_1_impl_parent_implementedSystem_port_1_cast);

SharedReg290_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg290_out;
SharedReg366_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg366_out;
SharedReg673_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg673_out;
SharedReg530_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg530_out;
SharedReg15_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg15_out;
SharedReg14_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg14_out;
SharedReg435_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg435_out;
SharedReg622_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg622_out;
SharedReg663_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg663_out;
Delay11No31_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_10_cast <= Delay11No31_out;
SharedReg529_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg529_out;
SharedReg674_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg674_out;
SharedReg622_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg622_out;
Delay16No1_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_14_cast <= Delay16No1_out;
   MUX_Add40_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg290_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg366_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg529_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg674_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg622_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay16No1_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg673_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg530_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg15_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg14_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg435_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg622_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg663_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay11No31_out_to_MUX_Add40_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add40_1_impl_0_out);

   Delay1No104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_1_impl_0_out,
                 Y => Delay1No104_out);

SharedReg673_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg673_out;
SharedReg475_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg475_out;
SharedReg663_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg663_out;
SharedReg673_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg673_out;
SharedReg31_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg31_out;
SharedReg30_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg30_out;
SharedReg454_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg454_out;
SharedReg663_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg663_out;
SharedReg398_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg398_out;
SharedReg291_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg291_out;
SharedReg621_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg621_out;
SharedReg289_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg289_out;
Delay15No36_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_13_cast <= Delay15No36_out;
SharedReg663_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg663_out;
   MUX_Add40_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg673_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg475_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg621_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg289_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay15No36_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg663_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg663_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg673_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg31_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg30_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg454_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg663_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg398_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg291_out_to_MUX_Add40_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add40_1_impl_1_out);

   Delay1No105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_1_impl_1_out,
                 Y => Delay1No105_out);

Delay1No106_out_to_Add40_2_impl_parent_implementedSystem_port_0_cast <= Delay1No106_out;
Delay1No107_out_to_Add40_2_impl_parent_implementedSystem_port_1_cast <= Delay1No107_out;
   Add40_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add40_2_impl_out,
                 X => Delay1No106_out_to_Add40_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No107_out_to_Add40_2_impl_parent_implementedSystem_port_1_cast);

SharedReg572_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg572_out;
SharedReg627_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg627_out;
Delay16No2_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_3_cast <= Delay16No2_out;
SharedReg572_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg572_out;
SharedReg369_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg369_out;
SharedReg571_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg571_out;
SharedReg600_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg600_out;
SharedReg15_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg15_out;
SharedReg14_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg14_out;
SharedReg439_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg439_out;
SharedReg600_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg600_out;
SharedReg665_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg665_out;
Delay11No32_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_13_cast <= Delay11No32_out;
SharedReg599_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg599_out;
   MUX_Add40_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg572_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg627_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg600_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg665_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay11No32_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg599_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => Delay16No2_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg572_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg369_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg571_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg600_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg15_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg14_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg439_out_to_MUX_Add40_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add40_2_impl_0_out);

   Delay1No106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_2_impl_0_out,
                 Y => Delay1No106_out);

SharedReg292_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg292_out;
Delay15No37_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_2_cast <= Delay15No37_out;
SharedReg627_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg627_out;
SharedReg664_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg664_out;
SharedReg534_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg534_out;
SharedReg665_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg665_out;
SharedReg571_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg571_out;
SharedReg31_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg31_out;
SharedReg30_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg30_out;
SharedReg457_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg457_out;
SharedReg627_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg627_out;
SharedReg402_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg402_out;
Delay3No252_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_13_cast <= Delay3No252_out;
SharedReg626_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg626_out;
   MUX_Add40_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg292_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay15No37_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg627_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg402_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay3No252_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg626_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg627_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg664_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg534_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg665_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg571_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg31_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg30_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg457_out_to_MUX_Add40_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add40_2_impl_1_out);

   Delay1No107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_2_impl_1_out,
                 Y => Delay1No107_out);

Delay1No108_out_to_Add40_3_impl_parent_implementedSystem_port_0_cast <= Delay1No108_out;
Delay1No109_out_to_Add40_3_impl_parent_implementedSystem_port_1_cast <= Delay1No109_out;
   Add40_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add40_3_impl_out,
                 X => Delay1No108_out_to_Add40_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No109_out_to_Add40_3_impl_parent_implementedSystem_port_1_cast);

SharedReg668_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg668_out;
Delay11No33_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_2_cast <= Delay11No33_out;
SharedReg538_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg538_out;
SharedReg668_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg668_out;
SharedReg606_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg606_out;
Delay16No3_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_6_cast <= Delay16No3_out;
SharedReg295_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg295_out;
SharedReg372_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg372_out;
SharedReg294_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg294_out;
SharedReg606_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg606_out;
SharedReg15_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg15_out;
SharedReg14_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg14_out;
SharedReg443_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg443_out;
SharedReg606_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg606_out;
   MUX_Add40_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg668_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay11No33_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg15_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg14_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg443_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg606_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg538_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg668_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg606_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay16No3_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg295_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg372_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg294_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg606_out_to_MUX_Add40_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add40_3_impl_0_out);

   Delay1No108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_3_impl_0_out,
                 Y => Delay1No108_out);

SharedReg405_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg405_out;
SharedReg302_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg302_out;
SharedReg605_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg605_out;
SharedReg294_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg294_out;
Delay15No38_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_5_cast <= Delay15No38_out;
SharedReg630_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg630_out;
SharedReg667_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg667_out;
SharedReg538_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg538_out;
SharedReg668_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg668_out;
SharedReg667_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg667_out;
SharedReg31_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg31_out;
SharedReg30_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg30_out;
SharedReg461_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg461_out;
SharedReg630_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg630_out;
   MUX_Add40_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg405_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg302_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg31_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg30_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg461_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg630_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg605_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg294_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay15No38_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg630_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg667_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg538_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg668_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg667_out_to_MUX_Add40_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add40_3_impl_1_out);

   Delay1No109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_3_impl_1_out,
                 Y => Delay1No109_out);

Delay1No110_out_to_Add40_4_impl_parent_implementedSystem_port_0_cast <= Delay1No110_out;
Delay1No111_out_to_Add40_4_impl_parent_implementedSystem_port_1_cast <= Delay1No111_out;
   Add40_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add40_4_impl_out,
                 X => Delay1No110_out_to_Add40_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No111_out_to_Add40_4_impl_parent_implementedSystem_port_1_cast);

SharedReg466_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg466_out;
SharedReg636_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg636_out;
SharedReg612_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg612_out;
Delay11No34_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_4_cast <= Delay11No34_out;
SharedReg486_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg486_out;
SharedReg636_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg636_out;
SharedReg612_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg612_out;
Delay16No4_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_8_cast <= Delay16No4_out;
SharedReg735_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg735_out;
SharedReg375_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg375_out;
SharedReg734_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg734_out;
SharedReg612_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg612_out;
SharedReg15_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg15_out;
SharedReg14_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg14_out;
   MUX_Add40_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg466_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg636_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg734_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg612_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg15_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg14_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg612_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay11No34_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg486_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg636_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg612_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay16No4_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg735_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg375_out_to_MUX_Add40_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add40_4_impl_0_out);

   Delay1No110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_4_impl_0_out,
                 Y => Delay1No110_out);

SharedReg486_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg486_out;
SharedReg677_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg677_out;
SharedReg428_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg428_out;
SharedReg678_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg678_out;
SharedReg542_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg542_out;
SharedReg734_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg734_out;
Delay15No39_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_7_cast <= Delay15No39_out;
SharedReg636_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg636_out;
SharedReg676_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg676_out;
SharedReg486_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg486_out;
SharedReg636_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg636_out;
SharedReg734_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg734_out;
SharedReg31_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg31_out;
SharedReg30_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg30_out;
   MUX_Add40_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg486_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg677_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg636_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg734_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg31_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg30_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg428_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg678_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg542_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg734_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay15No39_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg636_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg676_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg486_out_to_MUX_Add40_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Add40_4_impl_1_out);

   Delay1No111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add40_4_impl_1_out,
                 Y => Delay1No111_out);

Delay1No112_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast <= Delay1No112_out;
Delay1No113_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast <= Delay1No113_out;
   Product4_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_0_impl_out,
                 X => Delay1No112_out_to_Product4_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No113_out_to_Product4_0_impl_parent_implementedSystem_port_1_cast);

SharedReg849_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg849_out;
SharedReg792_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg792_out;
SharedReg787_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg787_out;
SharedReg63_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg63_out;
SharedReg812_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg812_out;
SharedReg798_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg798_out;
SharedReg821_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg821_out;
SharedReg777_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg777_out;
SharedReg778_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg778_out;
SharedReg492_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg492_out;
SharedReg62_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg62_out;
SharedReg783_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg783_out;
SharedReg784_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg784_out;
SharedReg790_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg790_out;
   MUX_Product4_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg849_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg792_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg62_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg783_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg784_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg790_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg787_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg63_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg812_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg798_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg821_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg777_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg778_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg492_out_to_MUX_Product4_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product4_0_impl_0_out);

   Delay1No112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_0_impl_0_out,
                 Y => Delay1No112_out);

SharedReg708_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg708_out;
SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg32_out;
Delay9No_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast <= Delay9No_out;
SharedReg811_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg811_out;
SharedReg34_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg34_out;
SharedReg66_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg66_out;
SharedReg679_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg679_out;
SharedReg63_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg63_out;
SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg33_out;
SharedReg829_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg829_out;
SharedReg805_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg805_out;
SharedReg63_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg63_out;
SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg33_out;
SharedReg62_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg62_out;
   MUX_Product4_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg708_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg32_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg805_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg63_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg62_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => Delay9No_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg811_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg34_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg66_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg679_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg63_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg33_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg829_out_to_MUX_Product4_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product4_0_impl_1_out);

   Delay1No113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_0_impl_1_out,
                 Y => Delay1No113_out);

Delay1No114_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast <= Delay1No114_out;
Delay1No115_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast <= Delay1No115_out;
   Product4_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_1_impl_out,
                 X => Delay1No114_out_to_Product4_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No115_out_to_Product4_1_impl_parent_implementedSystem_port_1_cast);

SharedReg804_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg804_out;
SharedReg637_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg637_out;
SharedReg843_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg843_out;
SharedReg679_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg679_out;
SharedReg817_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg817_out;
SharedReg787_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg787_out;
SharedReg862_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg862_out;
SharedReg575_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg575_out;
SharedReg239_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg239_out;
SharedReg779_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg779_out;
SharedReg803_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg803_out;
SharedReg778_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg778_out;
SharedReg499_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg499_out;
SharedReg68_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg68_out;
   MUX_Product4_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg804_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg637_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg803_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg778_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg499_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg68_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg843_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg679_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg817_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg787_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg862_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg575_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg239_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg779_out_to_MUX_Product4_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product4_1_impl_0_out);

   Delay1No114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_1_impl_0_out,
                 Y => Delay1No114_out);

SharedReg37_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg37_out;
SharedReg842_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg842_out;
SharedReg704_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg704_out;
SharedReg816_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg816_out;
SharedReg738_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg738_out;
Delay9No1_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast <= Delay9No1_out;
SharedReg574_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg574_out;
SharedReg863_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg863_out;
SharedReg801_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg801_out;
SharedReg240_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg240_out;
SharedReg159_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg159_out;
SharedReg39_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg39_out;
SharedReg829_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg829_out;
SharedReg805_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg805_out;
   MUX_Product4_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg37_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg842_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg159_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg39_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg829_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg805_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg704_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg816_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg738_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay9No1_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg574_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg863_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg801_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg240_out_to_MUX_Product4_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product4_1_impl_1_out);

   Delay1No115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_1_impl_1_out,
                 Y => Delay1No115_out);

Delay1No116_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast <= Delay1No116_out;
Delay1No117_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast <= Delay1No117_out;
   Product4_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_2_impl_out,
                 X => Delay1No116_out_to_Product4_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No117_out_to_Product4_2_impl_parent_implementedSystem_port_1_cast);

SharedReg778_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg778_out;
SharedReg506_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg506_out;
SharedReg74_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg74_out;
SharedReg804_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg804_out;
SharedReg642_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg642_out;
SharedReg790_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg790_out;
SharedReg684_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg684_out;
SharedReg817_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg817_out;
SharedReg787_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg787_out;
SharedReg862_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg862_out;
SharedReg580_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg580_out;
SharedReg798_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg798_out;
SharedReg821_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg821_out;
SharedReg777_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg777_out;
   MUX_Product4_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg778_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg506_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg580_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg798_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg821_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg777_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg74_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg804_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg642_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg790_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg684_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg817_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg787_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg862_out_to_MUX_Product4_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product4_2_impl_0_out);

   Delay1No116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_2_impl_0_out,
                 Y => Delay1No116_out);

SharedReg45_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg45_out;
SharedReg829_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg829_out;
SharedReg805_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg805_out;
SharedReg43_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg43_out;
SharedReg842_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg842_out;
SharedReg74_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg74_out;
SharedReg816_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg816_out;
SharedReg746_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg746_out;
Delay9No2_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast <= Delay9No2_out;
SharedReg579_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg579_out;
SharedReg863_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg863_out;
SharedReg78_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg78_out;
SharedReg689_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg689_out;
SharedReg75_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg75_out;
   MUX_Product4_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg45_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg829_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg863_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg78_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg689_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg75_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg805_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg43_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg842_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg74_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg816_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg746_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay9No2_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg579_out_to_MUX_Product4_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product4_2_impl_1_out);

   Delay1No117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_2_impl_1_out,
                 Y => Delay1No117_out);

Delay1No118_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast <= Delay1No118_out;
Delay1No119_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast <= Delay1No119_out;
   Product4_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_3_impl_out,
                 X => Delay1No118_out_to_Product4_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No119_out_to_Product4_3_impl_parent_implementedSystem_port_1_cast);

SharedReg798_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg798_out;
SharedReg821_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg821_out;
SharedReg777_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg777_out;
SharedReg778_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg778_out;
SharedReg513_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg513_out;
SharedReg782_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg782_out;
SharedReg804_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg804_out;
SharedReg647_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg647_out;
SharedReg790_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg790_out;
SharedReg689_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg689_out;
SharedReg817_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg817_out;
SharedReg85_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg85_out;
SharedReg81_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg81_out;
SharedReg812_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg812_out;
   MUX_Product4_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg798_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg821_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg817_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg85_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg81_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg812_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg777_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg778_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg513_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg782_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg804_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg647_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg790_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg689_out_to_MUX_Product4_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product4_3_impl_0_out);

   Delay1No118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_3_impl_0_out,
                 Y => Delay1No118_out);

SharedReg84_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg84_out;
SharedReg694_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg694_out;
SharedReg81_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg81_out;
SharedReg51_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg51_out;
SharedReg829_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg829_out;
SharedReg101_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg101_out;
SharedReg49_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg49_out;
SharedReg842_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg842_out;
SharedReg80_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg80_out;
SharedReg816_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg816_out;
SharedReg754_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg754_out;
SharedReg810_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg810_out;
SharedReg811_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg811_out;
SharedReg52_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg52_out;
   MUX_Product4_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg84_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg694_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg754_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg810_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg811_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg52_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg81_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg51_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg829_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg101_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg49_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg842_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg80_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg816_out_to_MUX_Product4_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product4_3_impl_1_out);

   Delay1No119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_3_impl_1_out,
                 Y => Delay1No119_out);

Delay1No120_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast <= Delay1No120_out;
Delay1No121_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast <= Delay1No121_out;
   Product4_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product4_4_impl_out,
                 X => Delay1No120_out_to_Product4_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No121_out_to_Product4_4_impl_parent_implementedSystem_port_1_cast);

SharedReg87_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg87_out;
SharedReg862_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg862_out;
SharedReg590_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg590_out;
SharedReg266_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg266_out;
SharedReg779_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg779_out;
SharedReg778_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg778_out;
SharedReg855_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg855_out;
SharedReg781_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg781_out;
SharedReg783_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg783_out;
SharedReg695_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg695_out;
SharedReg835_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg835_out;
SharedReg849_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg849_out;
SharedReg694_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg694_out;
SharedReg817_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg817_out;
   MUX_Product4_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg87_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg862_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg835_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg849_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg694_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg817_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg590_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg266_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg779_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg778_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg855_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg781_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg783_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg695_out_to_MUX_Product4_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product4_4_impl_0_out);

   Delay1No120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_4_impl_0_out,
                 Y => Delay1No120_out);

SharedReg811_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg811_out;
SharedReg589_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg589_out;
SharedReg863_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg863_out;
SharedReg801_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg801_out;
SharedReg267_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg267_out;
SharedReg57_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg57_out;
SharedReg724_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg724_out;
SharedReg53_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg53_out;
SharedReg87_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg87_out;
SharedReg841_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg841_out;
SharedReg652_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg652_out;
SharedReg732_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg732_out;
SharedReg816_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg816_out;
SharedReg762_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg762_out;
   MUX_Product4_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg811_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg589_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg652_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg732_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg816_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg762_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg863_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg801_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg267_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg57_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg724_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg53_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg87_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg841_out_to_MUX_Product4_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product4_4_impl_1_out);

   Delay1No121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product4_4_impl_1_out,
                 Y => Delay1No121_out);

Delay1No122_out_to_Product11_1_impl_parent_implementedSystem_port_0_cast <= Delay1No122_out;
Delay1No123_out_to_Product11_1_impl_parent_implementedSystem_port_1_cast <= Delay1No123_out;
   Product11_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_1_impl_out,
                 X => Delay1No122_out_to_Product11_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No123_out_to_Product11_1_impl_parent_implementedSystem_port_1_cast);

SharedReg783_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg783_out;
SharedReg784_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg784_out;
SharedReg790_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg790_out;
SharedReg849_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg849_out;
SharedReg792_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg792_out;
SharedReg73_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg73_out;
SharedReg69_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg69_out;
SharedReg812_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg812_out;
SharedReg798_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg798_out;
SharedReg821_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg821_out;
SharedReg777_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg777_out;
SharedReg801_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg801_out;
SharedReg828_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg828_out;
SharedReg782_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg782_out;
   MUX_Product11_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg783_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg784_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg777_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg801_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg828_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg782_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg790_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg849_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg792_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg73_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg69_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg812_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg798_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg821_out_to_MUX_Product11_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product11_1_impl_0_out);

   Delay1No122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_1_impl_0_out,
                 Y => Delay1No122_out);

SharedReg69_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg69_out;
SharedReg39_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg39_out;
SharedReg68_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg68_out;
SharedReg714_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg714_out;
SharedReg38_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg38_out;
SharedReg810_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg810_out;
SharedReg811_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg811_out;
SharedReg40_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg40_out;
SharedReg72_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg72_out;
SharedReg684_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg684_out;
SharedReg69_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg69_out;
SharedReg39_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg39_out;
SharedReg334_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg334_out;
SharedReg95_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg95_out;
   MUX_Product11_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg69_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg39_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg69_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg39_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg334_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg95_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg68_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg714_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg38_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg810_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg811_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg40_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg72_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg684_out_to_MUX_Product11_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product11_1_impl_1_out);

   Delay1No123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_1_impl_1_out,
                 Y => Delay1No123_out);

Delay1No124_out_to_Product11_4_impl_parent_implementedSystem_port_0_cast <= Delay1No124_out;
Delay1No125_out_to_Product11_4_impl_parent_implementedSystem_port_1_cast <= Delay1No125_out;
   Product11_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product11_4_impl_out,
                 X => Delay1No124_out_to_Product11_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No125_out_to_Product11_4_impl_parent_implementedSystem_port_1_cast);

SharedReg788_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg788_out;
SharedReg812_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg812_out;
SharedReg798_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg798_out;
SharedReg821_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg821_out;
SharedReg777_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg777_out;
SharedReg801_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg801_out;
SharedReg520_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg520_out;
SharedReg86_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg86_out;
SharedReg783_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg783_out;
SharedReg804_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg804_out;
SharedReg652_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg652_out;
SharedReg854_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg854_out;
SharedReg792_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg792_out;
SharedReg787_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg787_out;
   MUX_Product11_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg788_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg812_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg652_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg854_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg792_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg787_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg798_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg821_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg777_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg801_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg520_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg86_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg783_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg804_out_to_MUX_Product11_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product11_4_impl_0_out);

   Delay1No124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_4_impl_0_out,
                 Y => Delay1No124_out);

Delay10No4_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_1_cast <= Delay10No4_out;
SharedReg58_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg58_out;
SharedReg90_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg90_out;
SharedReg699_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg699_out;
SharedReg87_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg87_out;
SharedReg57_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg57_out;
SharedReg829_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg829_out;
SharedReg805_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg805_out;
SharedReg129_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg129_out;
SharedReg55_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg55_out;
SharedReg842_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg842_out;
SharedReg732_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg732_out;
SharedReg56_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg56_out;
Delay9No4_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_14_cast <= Delay9No4_out;
   MUX_Product11_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay10No4_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg58_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg842_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg732_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg56_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay9No4_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg90_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg699_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg87_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg57_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg829_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg805_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg129_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg55_out_to_MUX_Product11_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product11_4_impl_1_out);

   Delay1No125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product11_4_impl_1_out,
                 Y => Delay1No125_out);

Delay1No126_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast <= Delay1No126_out;
Delay1No127_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast <= Delay1No127_out;
   Product21_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_0_impl_out,
                 X => Delay1No126_out_to_Product21_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No127_out_to_Product21_0_impl_parent_implementedSystem_port_1_cast);

SharedReg854_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg854_out;
SharedReg786_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg786_out;
SharedReg67_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg67_out;
SharedReg788_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg788_out;
SharedReg789_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg789_out;
SharedReg796_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg796_out;
SharedReg848_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg848_out;
SharedReg63_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg63_out;
SharedReg801_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg801_out;
SharedReg828_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg828_out;
SharedReg782_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg782_out;
SharedReg783_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg783_out;
SharedReg807_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg807_out;
SharedReg813_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg813_out;
   MUX_Product21_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg854_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg786_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg782_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg783_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg807_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg813_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg67_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg788_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg789_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg796_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg848_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg63_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg801_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg828_out_to_MUX_Product21_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product21_0_impl_0_out);

   Delay1No126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_0_impl_0_out,
                 Y => Delay1No126_out);

SharedReg708_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg708_out;
SharedReg682_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg682_out;
SharedReg810_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg810_out;
Delay10No_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast <= Delay10No_out;
SharedReg34_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg34_out;
SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg32_out;
SharedReg704_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg704_out;
SharedReg800_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg800_out;
SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg33_out;
SharedReg327_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg327_out;
SharedReg92_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg92_out;
SharedReg109_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg109_out;
SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg33_out;
SharedReg62_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg62_out;
   MUX_Product21_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg708_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg682_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg92_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg109_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg62_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg810_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay10No_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg34_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg32_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg704_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg800_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg33_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg327_out_to_MUX_Product21_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product21_0_impl_1_out);

   Delay1No127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_0_impl_1_out,
                 Y => Delay1No127_out);

Delay1No128_out_to_Product21_2_impl_parent_implementedSystem_port_0_cast <= Delay1No128_out;
Delay1No129_out_to_Product21_2_impl_parent_implementedSystem_port_1_cast <= Delay1No129_out;
   Product21_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_2_impl_out,
                 X => Delay1No128_out_to_Product21_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No129_out_to_Product21_2_impl_parent_implementedSystem_port_1_cast);

SharedReg801_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg801_out;
SharedReg828_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg828_out;
SharedReg782_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg782_out;
SharedReg783_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg783_out;
SharedReg784_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg784_out;
SharedReg813_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg813_out;
SharedReg849_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg849_out;
SharedReg792_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg792_out;
SharedReg79_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg79_out;
SharedReg75_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg75_out;
SharedReg812_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg812_out;
SharedReg796_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg796_out;
SharedReg848_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg848_out;
SharedReg75_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg75_out;
   MUX_Product21_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg801_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg828_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg812_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg796_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg848_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg75_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg782_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg783_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg784_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg813_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg849_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg792_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg79_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg75_out_to_MUX_Product21_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product21_2_impl_0_out);

   Delay1No128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_2_impl_0_out,
                 Y => Delay1No128_out);

SharedReg45_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg45_out;
SharedReg341_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg341_out;
SharedReg98_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg98_out;
SharedReg75_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg75_out;
SharedReg45_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg45_out;
SharedReg74_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg74_out;
SharedReg720_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg720_out;
SharedReg44_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg44_out;
SharedReg810_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg810_out;
SharedReg811_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg811_out;
SharedReg46_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg46_out;
SharedReg44_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg44_out;
SharedReg716_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg716_out;
SharedReg800_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg800_out;
   MUX_Product21_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg45_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg341_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg46_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg44_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg716_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg800_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg98_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg75_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg45_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg74_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg720_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg44_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg810_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg811_out_to_MUX_Product21_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product21_2_impl_1_out);

   Delay1No129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_2_impl_1_out,
                 Y => Delay1No129_out);

Delay1No130_out_to_Product21_3_impl_parent_implementedSystem_port_0_cast <= Delay1No130_out;
Delay1No131_out_to_Product21_3_impl_parent_implementedSystem_port_1_cast <= Delay1No131_out;
   Product21_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product21_3_impl_out,
                 X => Delay1No130_out_to_Product21_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No131_out_to_Product21_3_impl_parent_implementedSystem_port_1_cast);

SharedReg796_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg796_out;
SharedReg848_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg848_out;
SharedReg81_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg81_out;
SharedReg801_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg801_out;
SharedReg828_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg828_out;
SharedReg782_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg782_out;
SharedReg783_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg783_out;
SharedReg784_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg784_out;
SharedReg813_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg813_out;
SharedReg849_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg849_out;
SharedReg792_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg792_out;
SharedReg787_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg787_out;
SharedReg788_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg788_out;
SharedReg789_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg789_out;
   MUX_Product21_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg796_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg848_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg792_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg787_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg788_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg789_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg81_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg801_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg828_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg782_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg783_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg784_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg813_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg849_out_to_MUX_Product21_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product21_3_impl_0_out);

   Delay1No130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_3_impl_0_out,
                 Y => Delay1No130_out);

SharedReg50_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg50_out;
SharedReg722_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg722_out;
SharedReg800_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg800_out;
SharedReg51_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg51_out;
SharedReg348_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg348_out;
SharedReg122_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg122_out;
SharedReg81_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg81_out;
SharedReg51_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg51_out;
SharedReg80_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg80_out;
SharedReg726_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg726_out;
SharedReg50_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg50_out;
SharedReg101_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg101_out;
Delay10No3_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_13_cast <= Delay10No3_out;
SharedReg52_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg52_out;
   MUX_Product21_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg50_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg722_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg50_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg101_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay10No3_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg52_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg800_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg51_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg348_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg122_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg81_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg51_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg80_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg726_out_to_MUX_Product21_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product21_3_impl_1_out);

   Delay1No131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product21_3_impl_1_out,
                 Y => Delay1No131_out);

Delay1No132_out_to_Product31_1_impl_parent_implementedSystem_port_0_cast <= Delay1No132_out;
Delay1No133_out_to_Product31_1_impl_parent_implementedSystem_port_1_cast <= Delay1No133_out;
   Product31_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_1_impl_out,
                 X => Delay1No132_out_to_Product31_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No133_out_to_Product31_1_impl_parent_implementedSystem_port_1_cast);

SharedReg783_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg783_out;
SharedReg807_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg807_out;
SharedReg813_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg813_out;
SharedReg854_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg854_out;
SharedReg786_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg786_out;
SharedReg787_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg787_out;
SharedReg788_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg788_out;
SharedReg789_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg789_out;
SharedReg796_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg796_out;
SharedReg848_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg848_out;
SharedReg69_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg69_out;
SharedReg830_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg830_out;
SharedReg828_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg828_out;
SharedReg782_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg782_out;
   MUX_Product31_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg783_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg807_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg69_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg830_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg828_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg782_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg813_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg854_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg786_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg787_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg788_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg789_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg796_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg848_out_to_MUX_Product31_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product31_1_impl_0_out);

   Delay1No132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_1_impl_0_out,
                 Y => Delay1No132_out);

SharedReg114_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg114_out;
SharedReg39_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg39_out;
SharedReg68_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg68_out;
SharedReg714_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg714_out;
SharedReg687_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg687_out;
SharedReg95_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg95_out;
Delay10No1_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_7_cast <= Delay10No1_out;
SharedReg40_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg40_out;
SharedReg38_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg38_out;
SharedReg710_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg710_out;
SharedReg800_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg800_out;
SharedReg552_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg552_out;
SharedReg499_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg499_out;
SharedReg112_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg112_out;
   MUX_Product31_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg114_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg39_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg800_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg552_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg499_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg112_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg68_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg714_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg687_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg95_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay10No1_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg40_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg38_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg710_out_to_MUX_Product31_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product31_1_impl_1_out);

   Delay1No133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_1_impl_1_out,
                 Y => Delay1No133_out);

Delay1No134_out_to_Product31_4_impl_parent_implementedSystem_port_0_cast <= Delay1No134_out;
Delay1No135_out_to_Product31_4_impl_parent_implementedSystem_port_1_cast <= Delay1No135_out;
   Product31_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product31_4_impl_out,
                 X => Delay1No134_out_to_Product31_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No135_out_to_Product31_4_impl_parent_implementedSystem_port_1_cast);

SharedReg788_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg788_out;
SharedReg789_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg789_out;
SharedReg796_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg796_out;
SharedReg848_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg848_out;
SharedReg87_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg87_out;
SharedReg830_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg830_out;
SharedReg828_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg828_out;
SharedReg782_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg782_out;
SharedReg129_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg129_out;
SharedReg784_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg784_out;
SharedReg790_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg790_out;
SharedReg808_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg808_out;
SharedReg786_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg786_out;
SharedReg91_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg91_out;
   MUX_Product31_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg788_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg789_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg790_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg808_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg786_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg91_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg796_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg848_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg87_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg830_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg828_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg782_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg129_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg784_out_to_MUX_Product31_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product31_4_impl_0_out);

   Delay1No134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_4_impl_0_out,
                 Y => Delay1No134_out);

SharedReg87_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg87_out;
SharedReg58_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg58_out;
SharedReg56_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg56_out;
SharedReg728_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg728_out;
SharedReg800_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg800_out;
SharedReg567_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg567_out;
SharedReg355_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg355_out;
SharedReg104_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg104_out;
SharedReg806_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg806_out;
SharedReg57_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg57_out;
SharedReg86_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg86_out;
SharedReg60_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg60_out;
SharedReg702_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg702_out;
SharedReg810_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg810_out;
   MUX_Product31_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg87_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg58_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg86_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg60_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg702_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg810_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg56_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg728_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg800_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg567_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg355_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg104_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg806_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg57_out_to_MUX_Product31_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product31_4_impl_1_out);

   Delay1No135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product31_4_impl_1_out,
                 Y => Delay1No135_out);

Delay1No136_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast <= Delay1No136_out;
Delay1No137_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast <= Delay1No137_out;
   Subtract2_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_0_impl_out,
                 X => Delay1No136_out_to_Subtract2_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No137_out_to_Subtract2_0_impl_parent_implementedSystem_port_1_cast);

SharedReg303_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg303_out;
SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg6_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg6_out;
SharedReg413_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg413_out;
SharedReg284_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg284_out;
SharedReg471_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg471_out;
SharedReg284_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg284_out;
SharedReg283_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg283_out;
SharedReg303_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg303_out;
SharedReg362_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg362_out;
SharedReg393_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg393_out;
SharedReg361_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg361_out;
SharedReg282_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg282_out;
SharedReg303_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg303_out;
   MUX_Subtract2_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg303_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg393_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg361_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg282_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg303_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg6_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg413_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg284_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg471_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg284_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg283_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg303_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg362_out_to_MUX_Subtract2_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract2_0_impl_0_out);

   Delay1No136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_0_out,
                 Y => Delay1No136_out);

SharedReg393_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg393_out;
SharedReg16_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg16_out;
SharedReg22_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg22_out;
SharedReg363_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg363_out;
Delay5No10_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast <= Delay5No10_out;
SharedReg619_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg619_out;
Delay10No25_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast <= Delay10No25_out;
SharedReg304_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg304_out;
SharedReg283_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg283_out;
SharedReg411_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg411_out;
SharedReg450_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg450_out;
SharedReg410_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg410_out;
SharedReg304_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg304_out;
SharedReg282_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg282_out;
   MUX_Subtract2_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg393_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg16_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg450_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg410_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg304_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg282_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg22_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg363_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay5No10_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg619_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay10No25_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg304_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg283_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg411_out_to_MUX_Subtract2_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract2_0_impl_1_out);

   Delay1No137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_0_impl_1_out,
                 Y => Delay1No137_out);

Delay1No138_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast <= Delay1No138_out;
Delay1No139_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast <= Delay1No139_out;
   Subtract2_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_1_impl_out,
                 X => Delay1No138_out_to_Subtract2_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No139_out_to_Subtract2_1_impl_parent_implementedSystem_port_1_cast);

SharedReg364_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg364_out;
SharedReg286_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg286_out;
SharedReg297_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg297_out;
SharedReg297_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg297_out;
SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg_out;
SharedReg6_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg6_out;
SharedReg399_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg399_out;
SharedReg299_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg299_out;
SharedReg476_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg476_out;
SharedReg299_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg299_out;
SharedReg287_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg287_out;
SharedReg317_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg317_out;
SharedReg365_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg365_out;
SharedReg396_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg396_out;
   MUX_Subtract2_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg364_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg286_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg287_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg317_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg365_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg396_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg297_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg297_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg6_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg399_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg299_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg476_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg299_out_to_MUX_Subtract2_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract2_1_impl_0_out);

   Delay1No138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_1_impl_0_out,
                 Y => Delay1No138_out);

SharedReg414_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg414_out;
SharedReg318_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg318_out;
SharedReg286_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg286_out;
SharedReg379_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg379_out;
SharedReg16_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg16_out;
SharedReg22_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg22_out;
SharedReg366_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg366_out;
Delay5No11_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast <= Delay5No11_out;
SharedReg624_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg624_out;
Delay10No26_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast <= Delay10No26_out;
SharedReg298_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg298_out;
SharedReg298_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg298_out;
SharedReg415_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg415_out;
SharedReg454_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg454_out;
   MUX_Subtract2_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg414_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg318_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg298_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg298_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg415_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg454_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg286_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg379_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg16_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg22_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg366_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay5No11_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg624_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay10No26_out_to_MUX_Subtract2_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract2_1_impl_1_out);

   Delay1No139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_1_impl_1_out,
                 Y => Delay1No139_out);

Delay1No140_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast <= Delay1No140_out;
Delay1No141_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast <= Delay1No141_out;
   Subtract2_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_2_impl_out,
                 X => Delay1No140_out_to_Subtract2_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No141_out_to_Subtract2_2_impl_parent_implementedSystem_port_1_cast);

SharedReg367_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg367_out;
SharedReg383_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg383_out;
SharedReg400_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg400_out;
SharedReg367_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg367_out;
SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg289_out;
SharedReg307_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg307_out;
SharedReg307_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg307_out;
SharedReg_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg_out;
SharedReg6_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg6_out;
SharedReg421_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg421_out;
SharedReg309_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg309_out;
SharedReg535_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg535_out;
SharedReg309_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg309_out;
SharedReg290_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg290_out;
   MUX_Subtract2_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg367_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg383_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg309_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg535_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg309_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg290_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg400_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg367_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg289_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg307_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg307_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg6_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg421_out_to_MUX_Subtract2_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract2_2_impl_0_out);

   Delay1No140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_2_impl_0_out,
                 Y => Delay1No140_out);

SharedReg308_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg308_out;
SharedReg440_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg440_out;
SharedReg457_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg457_out;
SharedReg418_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg418_out;
SharedReg308_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg308_out;
SharedReg289_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg289_out;
SharedReg400_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg400_out;
SharedReg16_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg16_out;
SharedReg22_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg22_out;
SharedReg384_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg384_out;
Delay5No12_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast <= Delay5No12_out;
Delay5No42_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast <= Delay5No42_out;
Delay10No27_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_13_cast <= Delay10No27_out;
SharedReg308_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg308_out;
   MUX_Subtract2_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg308_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg440_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay5No12_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay5No42_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay10No27_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg308_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg457_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg418_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg308_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg289_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg400_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg16_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg22_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg384_out_to_MUX_Subtract2_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract2_2_impl_1_out);

   Delay1No141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_2_impl_1_out,
                 Y => Delay1No141_out);

Delay1No142_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast <= Delay1No142_out;
Delay1No143_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast <= Delay1No143_out;
   Subtract2_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_3_impl_out,
                 X => Delay1No142_out_to_Subtract2_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No143_out_to_Subtract2_3_impl_parent_implementedSystem_port_1_cast);

SharedReg539_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg539_out;
SharedReg314_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg314_out;
SharedReg572_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg572_out;
SharedReg312_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg312_out;
SharedReg371_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg371_out;
SharedReg403_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg403_out;
SharedReg370_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg370_out;
SharedReg292_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg292_out;
SharedReg312_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg312_out;
SharedReg292_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg292_out;
SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg_out;
SharedReg6_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg6_out;
SharedReg406_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg406_out;
SharedReg314_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg314_out;
   MUX_Subtract2_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg539_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg314_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg6_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg406_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg314_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg572_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg312_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg371_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg403_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg370_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg292_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg312_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg292_out_to_MUX_Subtract2_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract2_3_impl_0_out);

   Delay1No142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_3_impl_0_out,
                 Y => Delay1No142_out);

Delay5No43_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast <= Delay5No43_out;
Delay10No28_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast <= Delay10No28_out;
SharedReg293_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg293_out;
SharedReg293_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg293_out;
SharedReg423_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg423_out;
SharedReg461_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg461_out;
SharedReg422_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg422_out;
SharedReg313_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg313_out;
SharedReg292_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg292_out;
SharedReg386_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg386_out;
SharedReg16_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg16_out;
SharedReg22_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg22_out;
SharedReg388_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg388_out;
Delay5No13_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_14_cast <= Delay5No13_out;
   MUX_Subtract2_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No43_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay10No28_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg16_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg22_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg388_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay5No13_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg293_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg293_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg423_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg461_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg422_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg313_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg292_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg386_out_to_MUX_Subtract2_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract2_3_impl_1_out);

   Delay1No143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_3_impl_1_out,
                 Y => Delay1No143_out);

Delay1No144_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast <= Delay1No144_out;
Delay1No145_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast <= Delay1No145_out;
   Subtract2_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract2_4_impl_out,
                 X => Delay1No144_out_to_Subtract2_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No145_out_to_Subtract2_4_impl_parent_implementedSystem_port_1_cast);

SharedReg429_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg429_out;
SharedReg323_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg323_out;
SharedReg467_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg467_out;
SharedReg296_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg296_out;
SharedReg301_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg301_out;
SharedReg321_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg321_out;
SharedReg374_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg374_out;
SharedReg407_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg407_out;
SharedReg373_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg373_out;
SharedReg294_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg294_out;
SharedReg321_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg321_out;
SharedReg321_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg321_out;
SharedReg_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg_out;
SharedReg6_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg6_out;
   MUX_Subtract2_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg429_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg323_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg321_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg321_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg6_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg467_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg296_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg301_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg321_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg374_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg407_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg373_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg294_out_to_MUX_Subtract2_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract2_4_impl_0_out);

   Delay1No144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_4_impl_0_out,
                 Y => Delay1No144_out);

SharedReg323_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg323_out;
Delay5No14_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast <= Delay5No14_out;
SharedReg545_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg545_out;
Delay10No29_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast <= Delay10No29_out;
SharedReg322_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg322_out;
SharedReg295_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg295_out;
SharedReg427_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg427_out;
SharedReg466_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg466_out;
SharedReg426_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg426_out;
SharedReg322_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg322_out;
SharedReg300_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg300_out;
SharedReg407_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg407_out;
SharedReg16_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg16_out;
SharedReg22_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg22_out;
   MUX_Subtract2_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg323_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay5No14_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg300_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg407_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg16_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg22_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg545_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay10No29_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg322_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg295_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg427_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg466_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg426_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg322_out_to_MUX_Subtract2_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract2_4_impl_1_out);

   Delay1No145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract2_4_impl_1_out,
                 Y => Delay1No145_out);

Delay1No146_out_to_Product5_0_impl_parent_implementedSystem_port_0_cast <= Delay1No146_out;
Delay1No147_out_to_Product5_0_impl_parent_implementedSystem_port_1_cast <= Delay1No147_out;
   Product5_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product5_0_impl_out,
                 X => Delay1No146_out_to_Product5_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No147_out_to_Product5_0_impl_parent_implementedSystem_port_1_cast);

SharedReg808_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg808_out;
SharedReg682_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg682_out;
SharedReg787_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg787_out;
SharedReg788_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg788_out;
SharedReg832_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg832_out;
SharedReg820_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg820_out;
SharedReg858_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg858_out;
SharedReg777_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg777_out;
SharedReg830_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg830_out;
SharedReg828_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg828_out;
SharedReg782_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg782_out;
SharedReg109_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg109_out;
SharedReg784_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg784_out;
SharedReg92_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg92_out;
   MUX_Product5_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg808_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg682_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg782_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg109_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg784_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg92_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg787_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg788_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg832_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg820_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg858_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg777_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg830_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg828_out_to_MUX_Product5_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product5_0_impl_0_out);

   Delay1No146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_0_impl_0_out,
                 Y => Delay1No146_out);

SharedReg36_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg36_out;
SharedReg809_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg809_out;
SharedReg92_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg92_out;
SharedReg63_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg63_out;
SharedReg640_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg640_out;
SharedReg66_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg66_out;
SharedReg736_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg736_out;
SharedReg93_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg93_out;
SharedReg547_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg547_out;
SharedReg492_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg492_out;
SharedReg107_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg107_out;
SharedReg806_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg806_out;
SharedReg134_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg134_out;
SharedReg813_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg813_out;
   MUX_Product5_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg36_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg809_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg107_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg806_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg134_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg813_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg92_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg63_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg640_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg66_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg736_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg93_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg547_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg492_out_to_MUX_Product5_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product5_0_impl_1_out);

   Delay1No147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_0_impl_1_out,
                 Y => Delay1No147_out);

Delay1No148_out_to_Product5_1_impl_parent_implementedSystem_port_0_cast <= Delay1No148_out;
Delay1No149_out_to_Product5_1_impl_parent_implementedSystem_port_1_cast <= Delay1No149_out;
   Product5_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product5_1_impl_out,
                 X => Delay1No148_out_to_Product5_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No149_out_to_Product5_1_impl_parent_implementedSystem_port_1_cast);

SharedReg114_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg114_out;
SharedReg784_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg784_out;
SharedReg95_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg95_out;
SharedReg808_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg808_out;
SharedReg687_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg687_out;
SharedReg787_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg787_out;
SharedReg788_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg788_out;
SharedReg832_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg832_out;
SharedReg820_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg820_out;
SharedReg858_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg858_out;
SharedReg777_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg777_out;
SharedReg830_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg830_out;
SharedReg829_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg829_out;
SharedReg805_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg805_out;
   MUX_Product5_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg114_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg784_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg777_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg830_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg829_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg805_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg95_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg808_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg687_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg787_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg788_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg832_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg820_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg858_out_to_MUX_Product5_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product5_1_impl_0_out);

   Delay1No148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_1_impl_0_out,
                 Y => Delay1No148_out);

SharedReg806_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg806_out;
SharedReg139_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg139_out;
SharedReg813_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg813_out;
SharedReg42_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg42_out;
SharedReg809_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg809_out;
SharedReg38_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg38_out;
SharedReg69_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg69_out;
SharedReg645_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg645_out;
SharedReg72_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg72_out;
SharedReg744_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg744_out;
SharedReg96_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg96_out;
SharedReg580_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg580_out;
SharedReg334_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg334_out;
SharedReg95_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg95_out;
   MUX_Product5_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg806_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg139_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg96_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg580_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg334_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg95_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg813_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg42_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg809_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg38_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg69_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg645_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg72_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg744_out_to_MUX_Product5_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product5_1_impl_1_out);

   Delay1No149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_1_impl_1_out,
                 Y => Delay1No149_out);

Delay1No150_out_to_Product5_2_impl_parent_implementedSystem_port_0_cast <= Delay1No150_out;
Delay1No151_out_to_Product5_2_impl_parent_implementedSystem_port_1_cast <= Delay1No151_out;
   Product5_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product5_2_impl_out,
                 X => Delay1No150_out_to_Product5_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No151_out_to_Product5_2_impl_parent_implementedSystem_port_1_cast);

SharedReg830_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg830_out;
SharedReg828_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg828_out;
SharedReg782_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg782_out;
SharedReg783_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg783_out;
SharedReg807_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg807_out;
SharedReg98_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg98_out;
SharedReg854_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg854_out;
SharedReg786_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg786_out;
SharedReg787_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg787_out;
SharedReg788_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg788_out;
SharedReg789_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg789_out;
SharedReg820_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg820_out;
SharedReg858_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg858_out;
SharedReg777_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg777_out;
   MUX_Product5_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg830_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg828_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg789_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg820_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg858_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg777_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg782_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg783_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg807_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg98_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg854_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg786_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg787_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg788_out_to_MUX_Product5_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product5_2_impl_0_out);

   Delay1No150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_2_impl_0_out,
                 Y => Delay1No150_out);

SharedReg557_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg557_out;
SharedReg506_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg506_out;
SharedReg117_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg117_out;
SharedReg119_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg119_out;
SharedReg45_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg45_out;
SharedReg813_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg813_out;
SharedReg720_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg720_out;
SharedReg692_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg692_out;
SharedReg98_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg98_out;
Delay10No2_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_10_cast <= Delay10No2_out;
SharedReg46_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg46_out;
SharedReg78_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg78_out;
SharedReg752_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg752_out;
SharedReg99_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg99_out;
   MUX_Product5_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg557_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg506_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg46_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg78_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg752_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg99_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg117_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg119_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg45_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg813_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg720_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg692_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg98_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay10No2_out_to_MUX_Product5_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product5_2_impl_1_out);

   Delay1No151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_2_impl_1_out,
                 Y => Delay1No151_out);

Delay1No152_out_to_Product5_3_impl_parent_implementedSystem_port_0_cast <= Delay1No152_out;
Delay1No153_out_to_Product5_3_impl_parent_implementedSystem_port_1_cast <= Delay1No153_out;
   Product5_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product5_3_impl_out,
                 X => Delay1No152_out_to_Product5_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No153_out_to_Product5_3_impl_parent_implementedSystem_port_1_cast);

SharedReg820_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg820_out;
SharedReg858_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg858_out;
SharedReg777_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg777_out;
SharedReg830_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg830_out;
SharedReg828_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg828_out;
SharedReg805_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg805_out;
SharedReg783_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg783_out;
SharedReg807_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg807_out;
SharedReg101_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg101_out;
SharedReg854_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg854_out;
SharedReg786_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg786_out;
SharedReg787_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg787_out;
SharedReg788_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg788_out;
SharedReg832_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg832_out;
   MUX_Product5_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg820_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg858_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg786_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg787_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg788_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg832_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg777_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg830_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg828_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg805_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg783_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg807_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg101_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg854_out_to_MUX_Product5_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product5_3_impl_0_out);

   Delay1No152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_3_impl_0_out,
                 Y => Delay1No152_out);

SharedReg84_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg84_out;
SharedReg760_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg760_out;
SharedReg102_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg102_out;
SharedReg562_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg562_out;
SharedReg513_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg513_out;
SharedReg101_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg101_out;
SharedReg124_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg124_out;
SharedReg51_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg51_out;
SharedReg813_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg813_out;
SharedReg726_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg726_out;
SharedReg697_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg697_out;
SharedReg50_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg50_out;
SharedReg81_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg81_out;
SharedReg655_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg655_out;
   MUX_Product5_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg84_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg760_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg697_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg50_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg81_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg655_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg102_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg562_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg513_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg101_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg124_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg51_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg813_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg726_out_to_MUX_Product5_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product5_3_impl_1_out);

   Delay1No153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_3_impl_1_out,
                 Y => Delay1No153_out);

Delay1No154_out_to_Product5_4_impl_parent_implementedSystem_port_0_cast <= Delay1No154_out;
Delay1No155_out_to_Product5_4_impl_parent_implementedSystem_port_1_cast <= Delay1No155_out;
   Product5_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product5_4_impl_out,
                 X => Delay1No154_out_to_Product5_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No155_out_to_Product5_4_impl_parent_implementedSystem_port_1_cast);

SharedReg794_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg794_out;
SharedReg832_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg832_out;
SharedReg820_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg820_out;
SharedReg858_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg858_out;
SharedReg777_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg777_out;
SharedReg830_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg830_out;
SharedReg828_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg828_out;
SharedReg782_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg782_out;
SharedReg824_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg824_out;
SharedReg807_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg807_out;
SharedReg813_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg813_out;
SharedReg785_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg785_out;
SharedReg702_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg702_out;
SharedReg787_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg787_out;
   MUX_Product5_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg794_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg832_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg813_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg785_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg702_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg787_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg820_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg858_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg777_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg830_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg828_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg782_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg824_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg807_out_to_MUX_Product5_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product5_4_impl_0_out);

   Delay1No154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_4_impl_0_out,
                 Y => Delay1No154_out);

SharedReg127_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg127_out;
SharedReg660_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg660_out;
SharedReg90_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg90_out;
SharedReg768_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg768_out;
SharedReg105_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg105_out;
SharedReg595_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg595_out;
SharedReg520_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg520_out;
SharedReg127_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg127_out;
SharedReg659_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg659_out;
SharedReg57_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg57_out;
SharedReg86_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg86_out;
SharedReg731_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg731_out;
SharedReg809_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg809_out;
SharedReg104_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg104_out;
   MUX_Product5_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg127_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg660_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg86_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg731_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg809_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg104_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg90_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg768_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg105_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg595_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg520_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg127_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg659_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg57_out_to_MUX_Product5_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product5_4_impl_1_out);

   Delay1No155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product5_4_impl_1_out,
                 Y => Delay1No155_out);

Delay1No156_out_to_Product12_0_impl_parent_implementedSystem_port_0_cast <= Delay1No156_out;
Delay1No157_out_to_Product12_0_impl_parent_implementedSystem_port_1_cast <= Delay1No157_out;
   Product12_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_0_impl_out,
                 X => Delay1No156_out_to_Product12_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No157_out_to_Product12_0_impl_parent_implementedSystem_port_1_cast);

SharedReg785_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg785_out;
SharedReg32_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg32_out;
SharedReg787_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg787_out;
SharedReg794_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg794_out;
SharedReg832_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg832_out;
SharedReg32_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg32_out;
SharedReg736_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg736_out;
SharedReg777_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg777_out;
SharedReg830_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg830_out;
SharedReg829_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg829_out;
SharedReg805_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg805_out;
SharedReg824_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg824_out;
SharedReg784_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg784_out;
SharedReg833_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg833_out;
   MUX_Product12_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg785_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg32_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg805_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg824_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg784_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg833_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg787_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg794_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg832_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg32_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg736_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg777_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg830_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg829_out_to_MUX_Product12_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product12_0_impl_0_out);

   Delay1No156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_0_impl_0_out,
                 Y => Delay1No156_out);

SharedReg707_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg707_out;
SharedReg814_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg814_out;
SharedReg32_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg32_out;
SharedReg107_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg107_out;
SharedReg576_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg576_out;
SharedReg818_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg818_out;
SharedReg860_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg860_out;
SharedReg108_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg108_out;
SharedReg575_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg575_out;
SharedReg327_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg327_out;
SharedReg92_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg92_out;
SharedReg639_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg639_out;
SharedReg159_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg159_out;
SharedReg637_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg637_out;
   MUX_Product12_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg707_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg814_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg92_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg639_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg159_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg637_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg32_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg107_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg576_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg818_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg860_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg108_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg575_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg327_out_to_MUX_Product12_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product12_0_impl_1_out);

   Delay1No157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_0_impl_1_out,
                 Y => Delay1No157_out);

Delay1No158_out_to_Product12_1_impl_parent_implementedSystem_port_0_cast <= Delay1No158_out;
Delay1No159_out_to_Product12_1_impl_parent_implementedSystem_port_1_cast <= Delay1No159_out;
   Product12_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_1_impl_out,
                 X => Delay1No158_out_to_Product12_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No159_out_to_Product12_1_impl_parent_implementedSystem_port_1_cast);

SharedReg824_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg824_out;
SharedReg784_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg784_out;
SharedReg833_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg833_out;
SharedReg785_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg785_out;
SharedReg38_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg38_out;
SharedReg810_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg810_out;
SharedReg794_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg794_out;
SharedReg832_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg832_out;
SharedReg38_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg38_out;
SharedReg744_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg744_out;
SharedReg777_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg777_out;
SharedReg837_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg837_out;
SharedReg845_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg845_out;
SharedReg112_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg112_out;
   MUX_Product12_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg824_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg784_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg777_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg837_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg845_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg112_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg833_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg785_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg38_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg810_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg794_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg832_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg38_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg744_out_to_MUX_Product12_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product12_1_impl_0_out);

   Delay1No158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_1_impl_0_out,
                 Y => Delay1No158_out);

SharedReg644_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg644_out;
SharedReg167_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg167_out;
SharedReg642_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg642_out;
SharedReg713_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg713_out;
SharedReg814_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg814_out;
SharedReg95_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg95_out;
SharedReg112_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg112_out;
SharedReg581_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg581_out;
SharedReg818_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg818_out;
SharedReg860_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg860_out;
SharedReg113_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg113_out;
SharedReg552_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg552_out;
SharedReg686_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg686_out;
SharedReg805_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg805_out;
   MUX_Product12_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg644_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg167_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg113_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg552_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg686_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg805_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg642_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg713_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg814_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg95_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg112_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg581_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg818_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg860_out_to_MUX_Product12_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product12_1_impl_1_out);

   Delay1No159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_1_impl_1_out,
                 Y => Delay1No159_out);

Delay1No160_out_to_Product12_2_impl_parent_implementedSystem_port_0_cast <= Delay1No160_out;
Delay1No161_out_to_Product12_2_impl_parent_implementedSystem_port_1_cast <= Delay1No161_out;
   Product12_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_2_impl_out,
                 X => Delay1No160_out_to_Product12_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No161_out_to_Product12_2_impl_parent_implementedSystem_port_1_cast);

SharedReg830_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg830_out;
SharedReg829_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg829_out;
SharedReg805_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg805_out;
SharedReg119_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg119_out;
SharedReg784_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg784_out;
SharedReg833_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg833_out;
SharedReg808_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg808_out;
SharedReg692_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg692_out;
SharedReg787_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg787_out;
SharedReg788_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg788_out;
SharedReg832_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg832_out;
SharedReg44_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg44_out;
SharedReg752_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg752_out;
SharedReg777_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg777_out;
   MUX_Product12_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg830_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg829_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg832_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg44_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg752_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg777_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg805_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg119_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg784_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg833_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg808_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg692_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg787_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg788_out_to_MUX_Product12_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product12_2_impl_0_out);

   Delay1No160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_2_impl_0_out,
                 Y => Delay1No160_out);

SharedReg585_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg585_out;
SharedReg341_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg341_out;
SharedReg98_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg98_out;
SharedReg806_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg806_out;
SharedReg144_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg144_out;
SharedReg647_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg647_out;
SharedReg48_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg48_out;
SharedReg809_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg809_out;
SharedReg44_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg44_out;
SharedReg75_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg75_out;
SharedReg650_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg650_out;
SharedReg818_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg818_out;
SharedReg860_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg860_out;
SharedReg118_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg118_out;
   MUX_Product12_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg585_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg341_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg650_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg818_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg860_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg118_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg98_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg806_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg144_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg647_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg48_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg809_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg44_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg75_out_to_MUX_Product12_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product12_2_impl_1_out);

   Delay1No161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_2_impl_1_out,
                 Y => Delay1No161_out);

Delay1No162_out_to_Product12_3_impl_parent_implementedSystem_port_0_cast <= Delay1No162_out;
Delay1No163_out_to_Product12_3_impl_parent_implementedSystem_port_1_cast <= Delay1No163_out;
   Product12_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_3_impl_out,
                 X => Delay1No162_out_to_Product12_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No163_out_to_Product12_3_impl_parent_implementedSystem_port_1_cast);

SharedReg50_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg50_out;
SharedReg760_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg760_out;
SharedReg777_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg777_out;
SharedReg830_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg830_out;
SharedReg829_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg829_out;
SharedReg122_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg122_out;
SharedReg124_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg124_out;
SharedReg784_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg784_out;
SharedReg833_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg833_out;
SharedReg808_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg808_out;
SharedReg697_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg697_out;
SharedReg810_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg810_out;
SharedReg794_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg794_out;
SharedReg832_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg832_out;
   MUX_Product12_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg50_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg760_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg697_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg810_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg794_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg832_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg777_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg830_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg829_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg122_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg124_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg784_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg833_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg808_out_to_MUX_Product12_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product12_3_impl_0_out);

   Delay1No162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_3_impl_0_out,
                 Y => Delay1No162_out);

SharedReg818_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg818_out;
SharedReg860_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg860_out;
SharedReg123_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg123_out;
SharedReg590_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg590_out;
SharedReg348_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg348_out;
SharedReg805_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg805_out;
SharedReg806_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg806_out;
SharedReg149_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg149_out;
SharedReg652_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg652_out;
SharedReg54_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg54_out;
SharedReg809_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg809_out;
SharedReg101_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg101_out;
SharedReg122_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg122_out;
SharedReg591_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg591_out;
   MUX_Product12_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg818_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg860_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg809_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg101_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg122_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg591_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg123_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg590_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg348_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg805_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg806_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg149_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg652_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg54_out_to_MUX_Product12_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product12_3_impl_1_out);

   Delay1No163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_3_impl_1_out,
                 Y => Delay1No163_out);

Delay1No164_out_to_Product12_4_impl_parent_implementedSystem_port_0_cast <= Delay1No164_out;
Delay1No165_out_to_Product12_4_impl_parent_implementedSystem_port_1_cast <= Delay1No165_out;
   Product12_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product12_4_impl_out,
                 X => Delay1No164_out_to_Product12_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No165_out_to_Product12_4_impl_parent_implementedSystem_port_1_cast);

SharedReg127_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg127_out;
SharedReg832_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg832_out;
SharedReg56_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg56_out;
SharedReg768_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg768_out;
SharedReg777_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg777_out;
SharedReg837_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg837_out;
SharedReg829_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg829_out;
SharedReg805_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg805_out;
SharedReg824_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg824_out;
SharedReg784_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg784_out;
SharedReg104_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg104_out;
SharedReg808_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg808_out;
SharedReg56_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg56_out;
SharedReg787_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg787_out;
   MUX_Product12_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg127_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg832_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg104_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg808_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg56_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg787_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg56_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg768_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg777_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg837_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg829_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg805_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg824_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg784_out_to_MUX_Product12_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product12_4_impl_0_out);

   Delay1No164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_4_impl_0_out,
                 Y => Delay1No164_out);

SharedReg816_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg816_out;
SharedReg596_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg596_out;
SharedReg818_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg818_out;
SharedReg860_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg860_out;
SharedReg128_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg128_out;
SharedReg567_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg567_out;
SharedReg355_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg355_out;
SharedReg104_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg104_out;
SharedReg701_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg701_out;
SharedReg154_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg154_out;
SharedReg813_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg813_out;
SharedReg731_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg731_out;
SharedReg814_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg814_out;
SharedReg56_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg56_out;
   MUX_Product12_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg816_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg596_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg813_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg731_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg814_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg56_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg818_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg860_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg128_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg567_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg355_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg104_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg701_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg154_out_to_MUX_Product12_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product12_4_impl_1_out);

   Delay1No165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product12_4_impl_1_out,
                 Y => Delay1No165_out);

Delay1No166_out_to_Product22_0_impl_parent_implementedSystem_port_0_cast <= Delay1No166_out;
Delay1No167_out_to_Product22_0_impl_parent_implementedSystem_port_1_cast <= Delay1No167_out;
   Product22_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_0_impl_out,
                 X => Delay1No166_out_to_Product22_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No167_out_to_Product22_0_impl_parent_implementedSystem_port_1_cast);

SharedReg808_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg808_out;
SharedReg792_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg792_out;
SharedReg810_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg810_out;
SharedReg107_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg107_out;
SharedReg839_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg839_out;
SharedReg796_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg796_out;
SharedReg776_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg776_out;
SharedReg800_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg800_out;
SharedReg837_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg837_out;
SharedReg845_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg845_out;
SharedReg107_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg107_out;
SharedReg824_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg824_out;
SharedReg807_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg807_out;
SharedReg840_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg840_out;
   MUX_Product22_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg808_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg792_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg107_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg824_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg807_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg840_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg810_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg107_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg839_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg796_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg776_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg800_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg837_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg845_out_to_MUX_Product22_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product22_0_impl_0_out);

   Delay1No166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_0_impl_0_out,
                 Y => Delay1No166_out);

SharedReg707_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg707_out;
SharedReg62_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg92_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg92_out;
SharedReg816_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg816_out;
SharedReg640_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg640_out;
SharedReg62_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg62_out;
SharedReg132_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg132_out;
SharedReg93_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg93_out;
SharedReg547_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg547_out;
SharedReg681_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg681_out;
SharedReg805_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg805_out;
SharedReg681_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg681_out;
SharedReg134_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg134_out;
SharedReg637_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg637_out;
   MUX_Product22_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg707_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg805_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg681_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg134_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg637_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg92_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg816_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg640_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg62_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg132_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg93_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg547_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg681_out_to_MUX_Product22_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product22_0_impl_1_out);

   Delay1No167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_0_impl_1_out,
                 Y => Delay1No167_out);

Delay1No168_out_to_Product22_1_impl_parent_implementedSystem_port_0_cast <= Delay1No168_out;
Delay1No169_out_to_Product22_1_impl_parent_implementedSystem_port_1_cast <= Delay1No169_out;
   Product22_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_1_impl_out,
                 X => Delay1No168_out_to_Product22_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No169_out_to_Product22_1_impl_parent_implementedSystem_port_1_cast);

SharedReg824_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg824_out;
SharedReg807_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg807_out;
SharedReg840_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg840_out;
SharedReg808_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg808_out;
SharedReg792_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg792_out;
SharedReg38_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg38_out;
SharedReg112_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg112_out;
SharedReg839_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg839_out;
SharedReg796_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg796_out;
SharedReg776_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg776_out;
SharedReg800_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg800_out;
SharedReg580_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg580_out;
SharedReg686_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg686_out;
SharedReg782_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg782_out;
   MUX_Product22_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg824_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg807_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg800_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg580_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg686_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg782_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg840_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg808_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg792_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg38_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg112_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg839_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg796_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg776_out_to_MUX_Product22_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product22_1_impl_0_out);

   Delay1No168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_1_impl_0_out,
                 Y => Delay1No168_out);

SharedReg686_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg686_out;
SharedReg139_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg139_out;
SharedReg642_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg642_out;
SharedReg713_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg713_out;
SharedReg68_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg68_out;
SharedReg810_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg810_out;
SharedReg816_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg816_out;
SharedReg645_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg645_out;
SharedReg68_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg68_out;
SharedReg137_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg137_out;
SharedReg96_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg96_out;
SharedReg837_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg837_out;
SharedReg847_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg847_out;
SharedReg96_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg96_out;
   MUX_Product22_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg686_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg139_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg96_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg837_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg847_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg96_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg642_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg713_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg68_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg810_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg816_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg645_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg68_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg137_out_to_MUX_Product22_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product22_1_impl_1_out);

   Delay1No169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_1_impl_1_out,
                 Y => Delay1No169_out);

Delay1No170_out_to_Product22_2_impl_parent_implementedSystem_port_0_cast <= Delay1No170_out;
Delay1No171_out_to_Product22_2_impl_parent_implementedSystem_port_1_cast <= Delay1No171_out;
   Product22_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_2_impl_out,
                 X => Delay1No170_out_to_Product22_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No171_out_to_Product22_2_impl_parent_implementedSystem_port_1_cast);

SharedReg837_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg837_out;
SharedReg845_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg845_out;
SharedReg117_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg117_out;
SharedReg824_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg824_out;
SharedReg784_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg784_out;
SharedReg840_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg840_out;
SharedReg785_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg785_out;
SharedReg44_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg44_out;
SharedReg810_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg810_out;
SharedReg794_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg794_out;
SharedReg832_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg832_out;
SharedReg796_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg796_out;
SharedReg776_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg776_out;
SharedReg800_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg800_out;
   MUX_Product22_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg837_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg845_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg832_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg796_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg776_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg800_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg117_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg824_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg784_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg840_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg785_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg44_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg810_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg794_out_to_MUX_Product22_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product22_2_impl_0_out);

   Delay1No170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_2_impl_0_out,
                 Y => Delay1No170_out);

SharedReg557_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg557_out;
SharedReg691_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg691_out;
SharedReg805_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg805_out;
SharedReg649_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg649_out;
SharedReg175_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg175_out;
SharedReg647_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg647_out;
SharedReg719_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg719_out;
SharedReg814_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg814_out;
SharedReg98_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg98_out;
SharedReg117_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg117_out;
SharedReg586_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg586_out;
SharedReg74_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg74_out;
SharedReg142_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg142_out;
SharedReg99_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg99_out;
   MUX_Product22_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg557_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg691_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg586_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg74_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg142_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg99_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg805_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg649_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg175_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg647_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg719_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg814_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg98_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg117_out_to_MUX_Product22_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product22_2_impl_1_out);

   Delay1No171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_2_impl_1_out,
                 Y => Delay1No171_out);

Delay1No172_out_to_Product22_3_impl_parent_implementedSystem_port_0_cast <= Delay1No172_out;
Delay1No173_out_to_Product22_3_impl_parent_implementedSystem_port_1_cast <= Delay1No173_out;
   Product22_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_3_impl_out,
                 X => Delay1No172_out_to_Product22_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No173_out_to_Product22_3_impl_parent_implementedSystem_port_1_cast);

SharedReg796_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg796_out;
SharedReg776_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg776_out;
SharedReg800_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg800_out;
SharedReg837_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg837_out;
SharedReg845_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg845_out;
SharedReg782_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg782_out;
SharedReg824_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg824_out;
SharedReg784_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg784_out;
SharedReg840_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg840_out;
SharedReg785_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg785_out;
SharedReg50_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg50_out;
SharedReg50_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg50_out;
SharedReg122_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg122_out;
SharedReg839_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg839_out;
   MUX_Product22_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg796_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg776_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg50_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg50_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg122_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg839_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg800_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg837_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg845_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg782_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg824_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg784_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg840_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg785_out_to_MUX_Product22_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product22_3_impl_0_out);

   Delay1No172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_3_impl_0_out,
                 Y => Delay1No172_out);

SharedReg80_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg80_out;
SharedReg147_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg147_out;
SharedReg102_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg102_out;
SharedReg562_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg562_out;
SharedReg696_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg696_out;
SharedReg102_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg102_out;
SharedReg654_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg654_out;
SharedReg183_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg183_out;
SharedReg652_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg652_out;
SharedReg725_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg725_out;
SharedReg814_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg814_out;
SharedReg810_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg810_out;
SharedReg816_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg816_out;
SharedReg655_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg655_out;
   MUX_Product22_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg80_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg147_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg814_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg810_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg816_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg655_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg102_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg562_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg696_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg102_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg654_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg183_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg652_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg725_out_to_MUX_Product22_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product22_3_impl_1_out);

   Delay1No173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_3_impl_1_out,
                 Y => Delay1No173_out);

Delay1No174_out_to_Product22_4_impl_parent_implementedSystem_port_0_cast <= Delay1No174_out;
Delay1No175_out_to_Product22_4_impl_parent_implementedSystem_port_1_cast <= Delay1No175_out;
   Product22_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product22_4_impl_out,
                 X => Delay1No174_out_to_Product22_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No175_out_to_Product22_4_impl_parent_implementedSystem_port_1_cast);

SharedReg794_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg794_out;
SharedReg839_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg839_out;
SharedReg796_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg796_out;
SharedReg776_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg776_out;
SharedReg800_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg800_out;
SharedReg595_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg595_out;
SharedReg845_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg845_out;
SharedReg127_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg127_out;
SharedReg827_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg827_out;
SharedReg784_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg784_out;
SharedReg833_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg833_out;
SharedReg785_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg785_out;
SharedReg792_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg792_out;
SharedReg810_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg810_out;
   MUX_Product22_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg794_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg839_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg833_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg785_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg792_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg810_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg796_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg776_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg800_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg595_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg845_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg127_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg827_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg784_out_to_MUX_Product22_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product22_4_impl_0_out);

   Delay1No174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_4_impl_0_out,
                 Y => Delay1No174_out);

SharedReg56_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg56_out;
SharedReg660_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg660_out;
SharedReg86_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg86_out;
SharedReg152_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg152_out;
SharedReg105_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg105_out;
SharedReg837_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg837_out;
SharedReg701_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg701_out;
SharedReg805_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg805_out;
SharedReg659_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg659_out;
SharedReg191_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg191_out;
SharedReg657_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg657_out;
SharedReg59_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg59_out;
SharedReg86_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg86_out;
SharedReg104_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg104_out;
   MUX_Product22_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg56_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg660_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg657_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg59_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg86_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg104_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg86_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg152_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg105_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg837_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg701_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg805_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg659_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg191_out_to_MUX_Product22_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product22_4_impl_1_out);

   Delay1No175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product22_4_impl_1_out,
                 Y => Delay1No175_out);

Delay1No176_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast <= Delay1No176_out;
Delay1No177_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast <= Delay1No177_out;
   Product32_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_0_impl_out,
                 X => Delay1No176_out_to_Product32_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No177_out_to_Product32_0_impl_parent_implementedSystem_port_1_cast);

SharedReg785_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg785_out;
SharedReg792_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg792_out;
SharedReg32_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg32_out;
SharedReg794_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg794_out;
SharedReg576_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg576_out;
SharedReg818_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg818_out;
SharedReg776_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg776_out;
SharedReg108_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg108_out;
SharedReg575_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg575_out;
SharedReg681_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg681_out;
SharedReg782_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg782_out;
SharedReg827_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg827_out;
SharedReg159_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg159_out;
SharedReg790_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg790_out;
   MUX_Product32_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg785_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg792_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg782_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg827_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg159_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg790_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg32_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg794_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg576_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg818_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg776_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg108_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg575_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg681_out_to_MUX_Product32_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product32_0_impl_0_out);

   Delay1No176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_0_impl_0_out,
                 Y => Delay1No176_out);

SharedReg35_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg35_out;
SharedReg92_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg92_out;
SharedReg810_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg810_out;
SharedReg32_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg32_out;
SharedReg839_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg839_out;
SharedReg62_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg62_out;
SharedReg157_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg157_out;
SharedReg800_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg800_out;
SharedReg837_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg837_out;
SharedReg847_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg847_out;
SharedReg93_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg93_out;
SharedReg639_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg639_out;
SharedReg807_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg807_out;
SharedReg32_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg32_out;
   MUX_Product32_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg35_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg92_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg93_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg639_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg807_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg32_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg810_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg32_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg839_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg62_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg157_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg800_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg837_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg847_out_to_MUX_Product32_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product32_0_impl_1_out);

   Delay1No177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_0_impl_1_out,
                 Y => Delay1No177_out);

Delay1No178_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast <= Delay1No178_out;
Delay1No179_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast <= Delay1No179_out;
   Product32_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_1_impl_out,
                 X => Delay1No178_out_to_Product32_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No179_out_to_Product32_1_impl_parent_implementedSystem_port_1_cast);

SharedReg827_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg827_out;
SharedReg167_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg167_out;
SharedReg790_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg790_out;
SharedReg785_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg785_out;
SharedReg792_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg792_out;
SharedReg793_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg793_out;
SharedReg794_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg794_out;
SharedReg581_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg581_out;
SharedReg818_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg818_out;
SharedReg776_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg776_out;
SharedReg113_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg113_out;
SharedReg844_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg844_out;
SharedReg779_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg779_out;
SharedReg805_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg805_out;
   MUX_Product32_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg827_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg167_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg113_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg844_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg779_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg805_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg790_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg785_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg792_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg793_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg794_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg581_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg818_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg776_out_to_MUX_Product32_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product32_1_impl_0_out);

   Delay1No178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_1_impl_0_out,
                 Y => Delay1No178_out);

SharedReg644_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg644_out;
SharedReg807_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg807_out;
SharedReg38_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg38_out;
SharedReg41_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg41_out;
SharedReg95_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg95_out;
SharedReg112_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg112_out;
SharedReg38_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg38_out;
SharedReg839_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg839_out;
SharedReg68_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg68_out;
SharedReg165_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg165_out;
SharedReg800_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg800_out;
SharedReg643_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg643_out;
SharedReg70_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg70_out;
SharedReg96_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg96_out;
   MUX_Product32_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg644_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg807_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg800_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg643_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg70_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg96_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg38_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg41_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg95_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg112_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg38_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg839_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg68_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg165_out_to_MUX_Product32_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product32_1_impl_1_out);

   Delay1No179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_1_impl_1_out,
                 Y => Delay1No179_out);

Delay1No180_out_to_Product32_2_impl_parent_implementedSystem_port_0_cast <= Delay1No180_out;
Delay1No181_out_to_Product32_2_impl_parent_implementedSystem_port_1_cast <= Delay1No181_out;
   Product32_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_2_impl_out,
                 X => Delay1No180_out_to_Product32_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No181_out_to_Product32_2_impl_parent_implementedSystem_port_1_cast);

SharedReg585_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg585_out;
SharedReg691_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg691_out;
SharedReg782_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg782_out;
SharedReg824_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg824_out;
SharedReg807_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg807_out;
SharedReg790_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg790_out;
SharedReg808_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg808_out;
SharedReg792_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg792_out;
SharedReg44_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg44_out;
SharedReg117_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg117_out;
SharedReg839_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg839_out;
SharedReg818_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg818_out;
SharedReg776_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg776_out;
SharedReg118_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg118_out;
   MUX_Product32_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg585_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg691_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg839_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg818_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg776_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg118_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg782_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg824_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg807_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg790_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg808_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg792_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg44_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg117_out_to_MUX_Product32_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product32_2_impl_0_out);

   Delay1No180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_2_impl_0_out,
                 Y => Delay1No180_out);

SharedReg837_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg837_out;
SharedReg847_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg847_out;
SharedReg99_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg99_out;
SharedReg691_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg691_out;
SharedReg144_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg144_out;
SharedReg44_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg44_out;
SharedReg719_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg719_out;
SharedReg74_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg74_out;
SharedReg810_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg810_out;
SharedReg816_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg816_out;
SharedReg650_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg650_out;
SharedReg74_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg74_out;
SharedReg173_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg173_out;
SharedReg800_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg800_out;
   MUX_Product32_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg837_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg847_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg650_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg74_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg173_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg800_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg99_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg691_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg144_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg44_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg719_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg74_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg810_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg816_out_to_MUX_Product32_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product32_2_impl_1_out);

   Delay1No181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_2_impl_1_out,
                 Y => Delay1No181_out);

Delay1No182_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast <= Delay1No182_out;
Delay1No183_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast <= Delay1No183_out;
   Product32_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_3_impl_out,
                 X => Delay1No182_out_to_Product32_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No183_out_to_Product32_3_impl_parent_implementedSystem_port_1_cast);

SharedReg818_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg818_out;
SharedReg776_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg776_out;
SharedReg123_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg123_out;
SharedReg590_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg590_out;
SharedReg696_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg696_out;
SharedReg805_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg805_out;
SharedReg824_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg824_out;
SharedReg807_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg807_out;
SharedReg790_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg790_out;
SharedReg808_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg808_out;
SharedReg792_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg792_out;
SharedReg793_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg793_out;
SharedReg794_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg794_out;
SharedReg591_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg591_out;
   MUX_Product32_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg818_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg776_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg792_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg793_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg794_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg591_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg123_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg590_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg696_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg805_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg824_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg807_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg790_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg808_out_to_MUX_Product32_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product32_3_impl_0_out);

   Delay1No182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_3_impl_0_out,
                 Y => Delay1No182_out);

SharedReg80_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg80_out;
SharedReg181_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg181_out;
SharedReg800_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg800_out;
SharedReg837_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg837_out;
SharedReg847_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg847_out;
SharedReg102_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg102_out;
SharedReg696_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg696_out;
SharedReg149_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg149_out;
SharedReg50_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg50_out;
SharedReg725_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg725_out;
SharedReg80_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg80_out;
SharedReg122_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg122_out;
SharedReg50_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg50_out;
SharedReg839_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg839_out;
   MUX_Product32_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg80_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg181_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg80_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg122_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg50_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg839_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg800_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg837_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg847_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg102_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg696_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg149_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg50_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg725_out_to_MUX_Product32_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product32_3_impl_1_out);

   Delay1No183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_3_impl_1_out,
                 Y => Delay1No183_out);

Delay1No184_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast <= Delay1No184_out;
Delay1No185_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast <= Delay1No185_out;
   Product32_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product32_4_impl_out,
                 X => Delay1No184_out_to_Product32_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No185_out_to_Product32_4_impl_parent_implementedSystem_port_1_cast);

SharedReg794_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg794_out;
SharedReg596_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg596_out;
SharedReg818_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg818_out;
SharedReg776_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg776_out;
SharedReg128_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg128_out;
SharedReg844_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg844_out;
SharedReg701_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg701_out;
SharedReg782_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg782_out;
SharedReg701_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg701_out;
SharedReg807_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg807_out;
SharedReg840_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg840_out;
SharedReg808_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg808_out;
SharedReg792_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg792_out;
SharedReg56_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg56_out;
   MUX_Product32_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg794_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg596_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg840_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg808_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg792_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg56_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg818_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg776_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg128_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg844_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg701_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg782_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg701_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg807_out_to_MUX_Product32_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product32_4_impl_0_out);

   Delay1No184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_4_impl_0_out,
                 Y => Delay1No184_out);

SharedReg86_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg86_out;
SharedReg839_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg839_out;
SharedReg86_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg86_out;
SharedReg189_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg189_out;
SharedReg800_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg800_out;
SharedReg658_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg658_out;
SharedReg847_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg847_out;
SharedReg105_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg105_out;
SharedReg827_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg827_out;
SharedReg154_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg154_out;
SharedReg657_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg657_out;
SharedReg59_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg59_out;
SharedReg104_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg104_out;
SharedReg810_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg810_out;
   MUX_Product32_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg86_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg839_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg657_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg59_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg104_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg810_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg86_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg189_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg800_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg658_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg847_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg105_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg827_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg154_out_to_MUX_Product32_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product32_4_impl_1_out);

   Delay1No185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product32_4_impl_1_out,
                 Y => Delay1No185_out);

Delay1No186_out_to_Product6_0_impl_parent_implementedSystem_port_0_cast <= Delay1No186_out;
Delay1No187_out_to_Product6_0_impl_parent_implementedSystem_port_1_cast <= Delay1No187_out;
   Product6_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_0_impl_out,
                 X => Delay1No186_out_to_Product6_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No187_out_to_Product6_0_impl_parent_implementedSystem_port_1_cast);

SharedReg808_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg808_out;
SharedReg814_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg814_out;
SharedReg793_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg793_out;
SharedReg794_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg794_out;
SharedReg795_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg795_out;
SharedReg796_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg796_out;
SharedReg799_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg799_out;
SharedReg822_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg822_out;
SharedReg844_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg844_out;
SharedReg779_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg779_out;
SharedReg805_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg805_out;
SharedReg681_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg681_out;
SharedReg784_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg784_out;
SharedReg790_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg790_out;
   MUX_Product6_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg808_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg814_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg805_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg681_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg784_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg790_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg793_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg794_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg795_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg796_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg799_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg822_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg844_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg779_out_to_MUX_Product6_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product6_0_impl_0_out);

   Delay1No186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_0_impl_0_out,
                 Y => Delay1No186_out);

SharedReg35_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg35_out;
SharedReg62_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg62_out;
SharedReg107_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg107_out;
SharedReg62_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg62_out;
SharedReg93_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg93_out;
SharedReg679_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg679_out;
SharedReg132_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg132_out;
SharedReg638_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg638_out;
SharedReg638_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg638_out;
SharedReg64_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg64_out;
SharedReg93_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg93_out;
SharedReg827_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg827_out;
SharedReg740_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg740_out;
SharedReg107_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg107_out;
   MUX_Product6_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg35_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg62_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg93_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg827_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg740_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg107_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg107_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg62_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg93_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg679_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg132_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg638_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg638_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg64_out_to_MUX_Product6_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product6_0_impl_1_out);

   Delay1No187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_0_impl_1_out,
                 Y => Delay1No187_out);

Delay1No188_out_to_Product6_1_impl_parent_implementedSystem_port_0_cast <= Delay1No188_out;
Delay1No189_out_to_Product6_1_impl_parent_implementedSystem_port_1_cast <= Delay1No189_out;
   Product6_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_1_impl_out,
                 X => Delay1No188_out_to_Product6_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No189_out_to_Product6_1_impl_parent_implementedSystem_port_1_cast);

SharedReg686_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg686_out;
SharedReg784_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg784_out;
SharedReg790_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg790_out;
SharedReg808_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg808_out;
SharedReg814_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg814_out;
SharedReg815_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg815_out;
SharedReg794_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg794_out;
SharedReg795_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg795_out;
SharedReg796_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg796_out;
SharedReg799_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg799_out;
SharedReg822_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg822_out;
SharedReg846_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg846_out;
SharedReg779_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg779_out;
SharedReg823_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg823_out;
   MUX_Product6_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg686_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg784_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg822_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg846_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg779_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg823_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg790_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg808_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg814_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg815_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg794_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg795_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg796_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg799_out_to_MUX_Product6_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product6_1_impl_0_out);

   Delay1No188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_1_impl_0_out,
                 Y => Delay1No188_out);

SharedReg827_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg827_out;
SharedReg748_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg748_out;
SharedReg112_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg112_out;
SharedReg41_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg41_out;
SharedReg68_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg68_out;
SharedReg112_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg112_out;
SharedReg68_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg68_out;
SharedReg96_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg96_out;
SharedReg684_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg684_out;
SharedReg137_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg137_out;
SharedReg643_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg643_out;
SharedReg643_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg643_out;
SharedReg97_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg97_out;
SharedReg710_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg710_out;
   MUX_Product6_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg827_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg748_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg643_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg643_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg97_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg710_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg112_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg41_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg68_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg112_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg68_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg96_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg684_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg137_out_to_MUX_Product6_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product6_1_impl_1_out);

   Delay1No189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_1_impl_1_out,
                 Y => Delay1No189_out);

Delay1No190_out_to_Product6_2_impl_parent_implementedSystem_port_0_cast <= Delay1No190_out;
Delay1No191_out_to_Product6_2_impl_parent_implementedSystem_port_1_cast <= Delay1No191_out;
   Product6_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_2_impl_out,
                 X => Delay1No190_out_to_Product6_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No191_out_to_Product6_2_impl_parent_implementedSystem_port_1_cast);

SharedReg844_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg844_out;
SharedReg779_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg779_out;
SharedReg805_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg805_out;
SharedReg827_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg827_out;
SharedReg175_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg175_out;
SharedReg790_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg790_out;
SharedReg785_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg785_out;
SharedReg792_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg792_out;
SharedReg793_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg793_out;
SharedReg794_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg794_out;
SharedReg586_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg586_out;
SharedReg796_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg796_out;
SharedReg799_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg799_out;
SharedReg822_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg822_out;
   MUX_Product6_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg844_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg779_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg586_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg796_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg799_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg822_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg805_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg827_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg175_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg790_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg785_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg792_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg793_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg794_out_to_MUX_Product6_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product6_2_impl_0_out);

   Delay1No190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_2_impl_0_out,
                 Y => Delay1No190_out);

SharedReg648_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg648_out;
SharedReg76_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg76_out;
SharedReg99_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg99_out;
SharedReg649_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg649_out;
SharedReg807_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg807_out;
SharedReg117_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg117_out;
SharedReg47_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg47_out;
SharedReg98_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg98_out;
SharedReg117_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg117_out;
SharedReg44_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg44_out;
SharedReg839_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg839_out;
SharedReg689_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg689_out;
SharedReg142_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg142_out;
SharedReg648_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg648_out;
   MUX_Product6_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg648_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg76_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg839_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg689_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg142_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg648_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg99_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg649_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg807_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg117_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg47_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg98_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg117_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg44_out_to_MUX_Product6_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product6_2_impl_1_out);

   Delay1No191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_2_impl_1_out,
                 Y => Delay1No191_out);

Delay1No192_out_to_Product6_3_impl_parent_implementedSystem_port_0_cast <= Delay1No192_out;
Delay1No193_out_to_Product6_3_impl_parent_implementedSystem_port_1_cast <= Delay1No193_out;
   Product6_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_3_impl_out,
                 X => Delay1No192_out_to_Product6_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No193_out_to_Product6_3_impl_parent_implementedSystem_port_1_cast);

SharedReg796_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg796_out;
SharedReg799_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg799_out;
SharedReg822_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg822_out;
SharedReg844_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg844_out;
SharedReg779_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg779_out;
SharedReg823_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg823_out;
SharedReg827_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg827_out;
SharedReg183_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg183_out;
SharedReg790_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg790_out;
SharedReg785_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg785_out;
SharedReg792_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg792_out;
SharedReg815_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg815_out;
SharedReg794_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg794_out;
SharedReg795_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg795_out;
   MUX_Product6_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg796_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg799_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg792_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg815_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg794_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg795_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg822_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg844_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg779_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg823_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg827_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg183_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg790_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg785_out_to_MUX_Product6_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product6_3_impl_0_out);

   Delay1No192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_3_impl_0_out,
                 Y => Delay1No192_out);

SharedReg694_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg694_out;
SharedReg147_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg147_out;
SharedReg653_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg653_out;
SharedReg653_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg653_out;
SharedReg82_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg82_out;
SharedReg722_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg722_out;
SharedReg654_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg654_out;
SharedReg807_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg807_out;
SharedReg122_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg122_out;
SharedReg53_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg53_out;
SharedReg101_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg101_out;
SharedReg122_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg122_out;
SharedReg80_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg80_out;
SharedReg102_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg102_out;
   MUX_Product6_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg694_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg147_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg101_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg122_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg80_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg102_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg653_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg653_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg82_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg722_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg654_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg807_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg122_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg53_out_to_MUX_Product6_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product6_3_impl_1_out);

   Delay1No193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_3_impl_1_out,
                 Y => Delay1No193_out);

Delay1No194_out_to_Product6_4_impl_parent_implementedSystem_port_0_cast <= Delay1No194_out;
Delay1No195_out_to_Product6_4_impl_parent_implementedSystem_port_1_cast <= Delay1No195_out;
   Product6_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product6_4_impl_out,
                 X => Delay1No194_out_to_Product6_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No195_out_to_Product6_4_impl_parent_implementedSystem_port_1_cast);

SharedReg816_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg816_out;
SharedReg795_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg795_out;
SharedReg796_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg796_out;
SharedReg799_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg799_out;
SharedReg822_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg822_out;
SharedReg846_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg846_out;
SharedReg779_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg779_out;
SharedReg805_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg805_out;
SharedReg783_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg783_out;
SharedReg191_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg191_out;
SharedReg790_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg790_out;
SharedReg785_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg785_out;
SharedReg814_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg814_out;
SharedReg793_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg793_out;
   MUX_Product6_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg816_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg795_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg790_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg785_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg814_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg793_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg796_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg799_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg822_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg846_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg779_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg805_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg783_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg191_out_to_MUX_Product6_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product6_4_impl_0_out);

   Delay1No194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_4_impl_0_out,
                 Y => Delay1No194_out);

SharedReg56_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg56_out;
SharedReg105_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg105_out;
SharedReg699_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg699_out;
SharedReg152_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg152_out;
SharedReg658_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg658_out;
SharedReg658_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg658_out;
SharedReg88_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg88_out;
SharedReg105_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg105_out;
SharedReg88_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg88_out;
SharedReg807_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg807_out;
SharedReg56_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg56_out;
SharedReg660_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg660_out;
SharedReg86_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg86_out;
SharedReg127_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg127_out;
   MUX_Product6_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg56_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg105_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg56_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg660_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg86_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg127_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg699_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg152_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg658_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg658_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg88_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg105_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg88_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg807_out_to_MUX_Product6_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product6_4_impl_1_out);

   Delay1No195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product6_4_impl_1_out,
                 Y => Delay1No195_out);

Delay1No196_out_to_Product23_0_impl_parent_implementedSystem_port_0_cast <= Delay1No196_out;
Delay1No197_out_to_Product23_0_impl_parent_implementedSystem_port_1_cast <= Delay1No197_out;
   Product23_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_0_impl_out,
                 X => Delay1No196_out_to_Product23_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No197_out_to_Product23_0_impl_parent_implementedSystem_port_1_cast);

SharedReg785_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg785_out;
SharedReg92_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg92_out;
SharedReg815_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg815_out;
SharedReg816_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg816_out;
SharedReg817_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg817_out;
SharedReg818_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg818_out;
SharedReg157_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg157_out;
SharedReg825_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg825_out;
SharedReg846_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg846_out;
SharedReg779_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg779_out;
SharedReg823_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg823_out;
SharedReg783_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg783_out;
SharedReg740_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg740_out;
SharedReg813_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg813_out;
   MUX_Product23_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg785_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg92_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg823_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg783_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg740_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg813_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg815_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg816_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg817_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg818_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg157_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg825_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg846_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg779_out_to_MUX_Product23_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product23_0_impl_0_out);

   Delay1No196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_0_impl_0_out,
                 Y => Delay1No196_out);

SharedReg640_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg640_out;
SharedReg814_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg814_out;
SharedReg107_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg107_out;
SharedReg32_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg32_out;
SharedReg93_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg93_out;
SharedReg679_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg679_out;
SharedReg799_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg799_out;
SharedReg638_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg638_out;
SharedReg638_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg638_out;
SharedReg94_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg94_out;
SharedReg704_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg704_out;
SharedReg64_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg64_out;
SharedReg807_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg807_out;
SharedReg32_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg32_out;
   MUX_Product23_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg640_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg814_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg704_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg64_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg807_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg32_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg107_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg32_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg93_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg679_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg799_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg638_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg638_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg94_out_to_MUX_Product23_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product23_0_impl_1_out);

   Delay1No197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_0_impl_1_out,
                 Y => Delay1No197_out);

Delay1No198_out_to_Product23_1_impl_parent_implementedSystem_port_0_cast <= Delay1No198_out;
Delay1No199_out_to_Product23_1_impl_parent_implementedSystem_port_1_cast <= Delay1No199_out;
   Product23_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_1_impl_out,
                 X => Delay1No198_out_to_Product23_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No199_out_to_Product23_1_impl_parent_implementedSystem_port_1_cast);

SharedReg783_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg783_out;
SharedReg748_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg748_out;
SharedReg813_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg813_out;
SharedReg785_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg785_out;
SharedReg95_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg95_out;
SharedReg831_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg831_out;
SharedReg816_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg816_out;
SharedReg817_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg817_out;
SharedReg818_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg818_out;
SharedReg165_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg165_out;
SharedReg825_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg825_out;
SharedReg859_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg859_out;
SharedReg802_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg802_out;
SharedReg826_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg826_out;
   MUX_Product23_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg783_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg748_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg825_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg859_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg802_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg826_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg813_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg785_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg95_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg831_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg816_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg817_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg818_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg165_out_to_MUX_Product23_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product23_1_impl_0_out);

   Delay1No198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_1_impl_0_out,
                 Y => Delay1No198_out);

SharedReg70_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg70_out;
SharedReg807_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg807_out;
SharedReg38_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg38_out;
SharedReg645_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg645_out;
SharedReg814_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg814_out;
SharedReg642_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg642_out;
SharedReg38_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg38_out;
SharedReg96_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg96_out;
SharedReg684_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg684_out;
SharedReg799_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg799_out;
SharedReg643_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg643_out;
SharedReg745_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg745_out;
SharedReg70_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg70_out;
SharedReg710_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg710_out;
   MUX_Product23_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg70_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg807_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg643_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg745_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg70_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg710_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg38_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg645_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg814_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg642_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg38_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg96_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg684_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg799_out_to_MUX_Product23_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product23_1_impl_1_out);

   Delay1No199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_1_impl_1_out,
                 Y => Delay1No199_out);

Delay1No200_out_to_Product23_2_impl_parent_implementedSystem_port_0_cast <= Delay1No200_out;
Delay1No201_out_to_Product23_2_impl_parent_implementedSystem_port_1_cast <= Delay1No201_out;
   Product23_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_2_impl_out,
                 X => Delay1No200_out_to_Product23_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No201_out_to_Product23_2_impl_parent_implementedSystem_port_1_cast);

SharedReg846_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg846_out;
SharedReg779_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg779_out;
SharedReg823_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg823_out;
SharedReg691_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg691_out;
SharedReg784_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg784_out;
SharedReg813_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg813_out;
SharedReg808_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg808_out;
SharedReg814_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg814_out;
SharedReg815_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg815_out;
SharedReg794_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg794_out;
SharedReg795_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg795_out;
SharedReg818_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg818_out;
SharedReg173_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg173_out;
SharedReg825_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg825_out;
   MUX_Product23_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg846_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg779_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg795_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg818_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg173_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg825_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg823_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg691_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg784_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg813_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg808_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg814_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg815_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg794_out_to_MUX_Product23_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product23_2_impl_0_out);

   Delay1No200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_2_impl_0_out,
                 Y => Delay1No200_out);

SharedReg648_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg648_out;
SharedReg100_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg100_out;
SharedReg716_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg716_out;
SharedReg827_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg827_out;
SharedReg756_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg756_out;
SharedReg44_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg44_out;
SharedReg47_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg47_out;
SharedReg74_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg74_out;
SharedReg117_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg117_out;
SharedReg74_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg74_out;
SharedReg99_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg99_out;
SharedReg689_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg689_out;
SharedReg799_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg799_out;
SharedReg648_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg648_out;
   MUX_Product23_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg648_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg100_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg99_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg689_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg799_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg648_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg716_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg827_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg756_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg44_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg47_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg74_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg117_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg74_out_to_MUX_Product23_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product23_2_impl_1_out);

   Delay1No201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_2_impl_1_out,
                 Y => Delay1No201_out);

Delay1No202_out_to_Product23_3_impl_parent_implementedSystem_port_0_cast <= Delay1No202_out;
Delay1No203_out_to_Product23_3_impl_parent_implementedSystem_port_1_cast <= Delay1No203_out;
   Product23_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_3_impl_out,
                 X => Delay1No202_out_to_Product23_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No203_out_to_Product23_3_impl_parent_implementedSystem_port_1_cast);

SharedReg818_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg818_out;
SharedReg181_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg181_out;
SharedReg825_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg825_out;
SharedReg846_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg846_out;
SharedReg779_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg779_out;
SharedReg826_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg826_out;
SharedReg696_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg696_out;
SharedReg784_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg784_out;
SharedReg813_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg813_out;
SharedReg808_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg808_out;
SharedReg814_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg814_out;
SharedReg831_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg831_out;
SharedReg816_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg816_out;
SharedReg817_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg817_out;
   MUX_Product23_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg818_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg181_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg814_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg831_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg816_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg817_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg825_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg846_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg779_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg826_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg696_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg784_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg813_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg808_out_to_MUX_Product23_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product23_3_impl_0_out);

   Delay1No202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_3_impl_0_out,
                 Y => Delay1No202_out);

SharedReg694_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg694_out;
SharedReg799_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg799_out;
SharedReg653_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg653_out;
SharedReg653_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg653_out;
SharedReg103_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg103_out;
SharedReg722_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg722_out;
SharedReg827_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg827_out;
SharedReg764_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg764_out;
SharedReg50_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg50_out;
SharedReg53_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg53_out;
SharedReg80_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg80_out;
SharedReg652_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg652_out;
SharedReg50_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg50_out;
SharedReg102_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg102_out;
   MUX_Product23_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg694_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg799_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg80_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg652_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg50_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg102_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg653_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg653_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg103_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg722_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg827_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg764_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg50_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg53_out_to_MUX_Product23_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product23_3_impl_1_out);

   Delay1No203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_3_impl_1_out,
                 Y => Delay1No203_out);

Delay1No204_out_to_Product23_4_impl_parent_implementedSystem_port_0_cast <= Delay1No204_out;
Delay1No205_out_to_Product23_4_impl_parent_implementedSystem_port_1_cast <= Delay1No205_out;
   Product23_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product23_4_impl_out,
                 X => Delay1No204_out_to_Product23_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No205_out_to_Product23_4_impl_parent_implementedSystem_port_1_cast);

SharedReg86_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg86_out;
SharedReg817_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg817_out;
SharedReg818_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg818_out;
SharedReg189_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg189_out;
SharedReg825_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg825_out;
SharedReg859_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg859_out;
SharedReg779_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg779_out;
SharedReg823_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg823_out;
SharedReg824_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg824_out;
SharedReg784_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg784_out;
SharedReg790_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg790_out;
SharedReg852_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg852_out;
SharedReg104_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg104_out;
SharedReg815_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg815_out;
   MUX_Product23_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg86_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg817_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg790_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg852_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg104_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg815_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg818_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg189_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg825_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg859_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg779_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg823_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg824_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg784_out_to_MUX_Product23_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product23_4_impl_0_out);

   Delay1No204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_4_impl_0_out,
                 Y => Delay1No204_out);

SharedReg816_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg816_out;
SharedReg105_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg105_out;
SharedReg699_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg699_out;
SharedReg799_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg799_out;
SharedReg658_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg658_out;
SharedReg769_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg769_out;
SharedReg106_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg106_out;
SharedReg728_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg728_out;
SharedReg769_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg769_out;
SharedReg772_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg772_out;
SharedReg127_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg127_out;
SharedReg597_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg597_out;
SharedReg814_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg814_out;
SharedReg127_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg127_out;
   MUX_Product23_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg816_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg105_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg127_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg597_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg814_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg127_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg699_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg799_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg658_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg769_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg106_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg728_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg769_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg772_out_to_MUX_Product23_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product23_4_impl_1_out);

   Delay1No205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product23_4_impl_1_out,
                 Y => Delay1No205_out);

Delay1No206_out_to_Product33_0_impl_parent_implementedSystem_port_0_cast <= Delay1No206_out;
Delay1No207_out_to_Product33_0_impl_parent_implementedSystem_port_1_cast <= Delay1No207_out;
   Product33_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_0_impl_out,
                 X => Delay1No206_out_to_Product33_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No207_out_to_Product33_0_impl_parent_implementedSystem_port_1_cast);

SharedReg852_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg852_out;
SharedReg835_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg835_out;
SharedReg831_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg831_out;
SharedReg62_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg62_out;
SharedReg797_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg797_out;
SharedReg742_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg742_out;
SharedReg776_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg776_out;
SharedReg680_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg680_out;
SharedReg859_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg859_out;
SharedReg802_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg802_out;
SharedReg826_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg826_out;
SharedReg824_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg824_out;
SharedReg65_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg65_out;
SharedReg107_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg107_out;
   MUX_Product33_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg852_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg835_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg826_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg824_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg65_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg107_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg831_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg62_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg797_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg742_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg776_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg680_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg859_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg802_out_to_MUX_Product33_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product33_0_impl_0_out);

   Delay1No206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_0_impl_0_out,
                 Y => Delay1No206_out);

SharedReg577_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg577_out;
SharedReg679_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg679_out;
SharedReg637_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg637_out;
SharedReg816_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg816_out;
SharedReg36_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg36_out;
SharedReg820_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg820_out;
SharedReg197_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg197_out;
SharedReg825_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg825_out;
SharedReg737_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg737_out;
SharedReg64_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg64_out;
SharedReg704_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg704_out;
SharedReg737_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg737_out;
SharedReg807_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg807_out;
SharedReg813_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg813_out;
   MUX_Product33_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg577_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg679_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg704_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg737_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg807_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg813_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg637_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg816_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg36_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg820_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg197_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg825_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg737_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg64_out_to_MUX_Product33_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product33_0_impl_1_out);

   Delay1No207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_0_impl_1_out,
                 Y => Delay1No207_out);

Delay1No208_out_to_Product33_1_impl_parent_implementedSystem_port_0_cast <= Delay1No208_out;
Delay1No209_out_to_Product33_1_impl_parent_implementedSystem_port_1_cast <= Delay1No209_out;
   Product33_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_1_impl_out,
                 X => Delay1No208_out_to_Product33_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No209_out_to_Product33_1_impl_parent_implementedSystem_port_1_cast);

SharedReg824_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg824_out;
SharedReg71_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg71_out;
SharedReg112_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg112_out;
SharedReg852_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg852_out;
SharedReg835_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg835_out;
SharedReg831_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg831_out;
SharedReg68_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg68_out;
SharedReg797_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg797_out;
SharedReg750_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg750_out;
SharedReg776_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg776_out;
SharedReg685_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg685_out;
SharedReg861_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg861_out;
SharedReg97_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg97_out;
SharedReg744_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg744_out;
   MUX_Product33_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg824_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg71_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg685_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg861_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg97_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg744_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg112_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg852_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg835_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg831_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg68_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg797_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg750_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg776_out_to_MUX_Product33_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product33_1_impl_0_out);

   Delay1No208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_1_impl_0_out,
                 Y => Delay1No208_out);

SharedReg745_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg745_out;
SharedReg807_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg807_out;
SharedReg813_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg813_out;
SharedReg582_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg582_out;
SharedReg684_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg684_out;
SharedReg684_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg684_out;
SharedReg816_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg816_out;
SharedReg42_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg42_out;
SharedReg820_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg820_out;
SharedReg205_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg205_out;
SharedReg825_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg825_out;
SharedReg745_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg745_out;
SharedReg802_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg802_out;
SharedReg826_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg826_out;
   MUX_Product33_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg745_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg807_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg825_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg745_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg802_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg826_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg813_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg582_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg684_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg684_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg816_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg42_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg820_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg205_out_to_MUX_Product33_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product33_1_impl_1_out);

   Delay1No209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_1_impl_1_out,
                 Y => Delay1No209_out);

Delay1No210_out_to_Product33_2_impl_parent_implementedSystem_port_0_cast <= Delay1No210_out;
Delay1No211_out_to_Product33_2_impl_parent_implementedSystem_port_1_cast <= Delay1No211_out;
   Product33_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_2_impl_out,
                 X => Delay1No210_out_to_Product33_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No211_out_to_Product33_2_impl_parent_implementedSystem_port_1_cast);

SharedReg859_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg859_out;
SharedReg802_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg802_out;
SharedReg826_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg826_out;
SharedReg783_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg783_out;
SharedReg756_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg756_out;
SharedReg117_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg117_out;
SharedReg785_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg785_out;
SharedReg98_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg98_out;
SharedReg831_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg831_out;
SharedReg816_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg816_out;
SharedReg817_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg817_out;
SharedReg758_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg758_out;
SharedReg776_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg776_out;
SharedReg690_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg690_out;
   MUX_Product33_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg859_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg802_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg817_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg758_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg776_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg690_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg826_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg783_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg756_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg117_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg785_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg98_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg831_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg816_out_to_MUX_Product33_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product33_2_impl_0_out);

   Delay1No210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_2_impl_0_out,
                 Y => Delay1No210_out);

SharedReg753_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg753_out;
SharedReg76_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg76_out;
SharedReg716_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg716_out;
SharedReg76_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg76_out;
SharedReg807_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg807_out;
SharedReg813_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg813_out;
SharedReg650_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg650_out;
SharedReg814_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg814_out;
SharedReg647_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg647_out;
SharedReg44_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg44_out;
SharedReg99_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg99_out;
SharedReg820_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg820_out;
SharedReg213_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg213_out;
SharedReg825_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg825_out;
   MUX_Product33_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg753_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg76_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg99_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg820_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg213_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg825_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg716_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg76_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg807_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg813_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg650_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg814_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg647_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg44_out_to_MUX_Product33_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product33_2_impl_1_out);

   Delay1No211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_2_impl_1_out,
                 Y => Delay1No211_out);

Delay1No212_out_to_Product33_3_impl_parent_implementedSystem_port_0_cast <= Delay1No212_out;
Delay1No213_out_to_Product33_3_impl_parent_implementedSystem_port_1_cast <= Delay1No213_out;
   Product33_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_3_impl_out,
                 X => Delay1No212_out_to_Product33_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No213_out_to_Product33_3_impl_parent_implementedSystem_port_1_cast);

SharedReg766_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg766_out;
SharedReg776_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg776_out;
SharedReg695_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg695_out;
SharedReg859_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg859_out;
SharedReg802_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg802_out;
SharedReg760_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg760_out;
SharedReg783_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg783_out;
SharedReg764_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg764_out;
SharedReg122_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg122_out;
SharedReg785_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg785_out;
SharedReg101_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg101_out;
SharedReg831_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg831_out;
SharedReg80_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg80_out;
SharedReg797_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg797_out;
   MUX_Product33_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg766_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg776_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg101_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg831_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg80_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg797_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg695_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg859_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg802_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg760_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg783_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg764_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg122_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg785_out_to_MUX_Product33_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product33_3_impl_0_out);

   Delay1No212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_3_impl_0_out,
                 Y => Delay1No212_out);

SharedReg820_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg820_out;
SharedReg221_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg221_out;
SharedReg825_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg825_out;
SharedReg761_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg761_out;
SharedReg82_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg82_out;
SharedReg826_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg826_out;
SharedReg82_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg82_out;
SharedReg807_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg807_out;
SharedReg813_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg813_out;
SharedReg655_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg655_out;
SharedReg814_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg814_out;
SharedReg694_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg694_out;
SharedReg816_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg816_out;
SharedReg54_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg54_out;
   MUX_Product33_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg820_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg221_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg814_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg694_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg816_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg54_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg825_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg761_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg82_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg826_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg82_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg807_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg813_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg655_out_to_MUX_Product33_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product33_3_impl_1_out);

   Delay1No213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_3_impl_1_out,
                 Y => Delay1No213_out);

Delay1No214_out_to_Product33_4_impl_parent_implementedSystem_port_0_cast <= Delay1No214_out;
Delay1No215_out_to_Product33_4_impl_parent_implementedSystem_port_1_cast <= Delay1No215_out;
   Product33_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product33_4_impl_out,
                 X => Delay1No214_out_to_Product33_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No215_out_to_Product33_4_impl_parent_implementedSystem_port_1_cast);

SharedReg794_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg794_out;
SharedReg797_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg797_out;
SharedReg774_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg774_out;
SharedReg776_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg776_out;
SharedReg700_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg700_out;
SharedReg861_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg861_out;
SharedReg802_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg802_out;
SharedReg826_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg826_out;
SharedReg850_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg850_out;
SharedReg772_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg772_out;
SharedReg813_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg813_out;
SharedReg857_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg857_out;
SharedReg835_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg835_out;
SharedReg831_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg831_out;
   MUX_Product33_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg794_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg797_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg813_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg857_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg835_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg831_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg774_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg776_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg700_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg861_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg802_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg826_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg850_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg772_out_to_MUX_Product33_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product33_4_impl_0_out);

   Delay1No214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_4_impl_0_out,
                 Y => Delay1No214_out);

SharedReg657_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg657_out;
SharedReg60_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg60_out;
SharedReg820_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg820_out;
SharedReg229_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg229_out;
SharedReg825_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg825_out;
SharedReg769_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg769_out;
SharedReg88_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg88_out;
SharedReg728_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg728_out;
SharedReg596_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg596_out;
SharedReg807_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg807_out;
SharedReg56_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg56_out;
SharedReg597_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg597_out;
SharedReg699_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg699_out;
SharedReg657_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg657_out;
   MUX_Product33_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg657_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg60_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg56_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg597_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg699_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg657_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg820_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg229_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg825_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg769_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg88_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg728_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg596_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg807_out_to_MUX_Product33_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product33_4_impl_1_out);

   Delay1No215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product33_4_impl_1_out,
                 Y => Delay1No215_out);

Delay1No216_out_to_Subtract4_0_impl_parent_implementedSystem_port_0_cast <= Delay1No216_out;
Delay1No217_out_to_Subtract4_0_impl_parent_implementedSystem_port_1_cast <= Delay1No217_out;
   Subtract4_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_0_impl_out,
                 X => Delay1No216_out_to_Subtract4_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No217_out_to_Subtract4_0_impl_parent_implementedSystem_port_1_cast);

SharedReg450_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg450_out;
SharedReg1_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1_out;
SharedReg7_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg7_out;
SharedReg362_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg362_out;
SharedReg283_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg283_out;
SharedReg393_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg393_out;
SharedReg361_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg361_out;
SharedReg452_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg452_out;
SharedReg632_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg632_out;
SharedReg282_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg282_out;
SharedReg526_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg526_out;
SharedReg430_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg430_out;
SharedReg361_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg361_out;
SharedReg431_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg431_out;
   MUX_Subtract4_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg450_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg526_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg430_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg361_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg431_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg7_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg362_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg283_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg393_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg361_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg452_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg632_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg282_out_to_MUX_Subtract4_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract4_0_impl_0_out);

   Delay1No216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_0_impl_0_out,
                 Y => Delay1No216_out);

SharedReg525_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg525_out;
SharedReg17_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg17_out;
SharedReg23_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg23_out;
SharedReg411_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg411_out;
SharedReg362_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg362_out;
SharedReg450_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg450_out;
SharedReg410_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg410_out;
SharedReg363_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg363_out;
SharedReg633_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg633_out;
Delay15No15_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_10_cast <= Delay15No15_out;
Delay16No5_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_11_cast <= Delay16No5_out;
SharedReg470_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg470_out;
SharedReg410_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg410_out;
SharedReg410_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg410_out;
   MUX_Subtract4_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg525_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg17_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay16No5_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg470_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg410_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg410_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg23_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg411_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg362_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg450_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg410_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg363_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg633_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay15No15_out_to_MUX_Subtract4_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract4_0_impl_1_out);

   Delay1No217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_0_impl_1_out,
                 Y => Delay1No217_out);

Delay1No218_out_to_Subtract4_1_impl_parent_implementedSystem_port_0_cast <= Delay1No218_out;
Delay1No219_out_to_Subtract4_1_impl_parent_implementedSystem_port_1_cast <= Delay1No219_out;
   Subtract4_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_1_impl_out,
                 X => Delay1No218_out_to_Subtract4_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No219_out_to_Subtract4_1_impl_parent_implementedSystem_port_1_cast);

SharedReg435_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg435_out;
SharedReg317_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg317_out;
SharedReg415_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg415_out;
SharedReg435_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg435_out;
SharedReg1_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1_out;
SharedReg7_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg7_out;
SharedReg365_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg365_out;
SharedReg298_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg298_out;
SharedReg396_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg396_out;
SharedReg317_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg317_out;
SharedReg455_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg455_out;
SharedReg662_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg662_out;
SharedReg297_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg297_out;
SharedReg530_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg530_out;
   MUX_Subtract4_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg435_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg317_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg455_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg662_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg297_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg530_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg415_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg435_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg7_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg365_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg298_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg396_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg317_out_to_MUX_Subtract4_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract4_1_impl_0_out);

   Delay1No218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_1_impl_0_out,
                 Y => Delay1No218_out);

SharedReg475_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg475_out;
SharedReg396_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg396_out;
SharedReg396_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg396_out;
SharedReg475_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg475_out;
SharedReg17_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg17_out;
SharedReg23_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg23_out;
SharedReg415_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg415_out;
SharedReg365_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg365_out;
SharedReg454_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg454_out;
SharedReg396_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg396_out;
SharedReg366_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg366_out;
SharedReg663_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg663_out;
Delay15No16_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_13_cast <= Delay15No16_out;
Delay16No6_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_14_cast <= Delay16No6_out;
   MUX_Subtract4_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg475_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg396_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg366_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg663_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay15No16_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => Delay16No6_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg396_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg475_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg17_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg23_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg415_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg365_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg454_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg396_out_to_MUX_Subtract4_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract4_1_impl_1_out);

   Delay1No219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_1_impl_1_out,
                 Y => Delay1No219_out);

Delay1No220_out_to_Subtract4_2_impl_parent_implementedSystem_port_0_cast <= Delay1No220_out;
Delay1No221_out_to_Subtract4_2_impl_parent_implementedSystem_port_1_cast <= Delay1No221_out;
   Subtract4_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_2_impl_out,
                 X => Delay1No220_out_to_Subtract4_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No221_out_to_Subtract4_2_impl_parent_implementedSystem_port_1_cast);

SharedReg664_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg664_out;
SharedReg289_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg289_out;
SharedReg535_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg535_out;
SharedReg439_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg439_out;
SharedReg367_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg367_out;
SharedReg440_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg440_out;
SharedReg457_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg457_out;
SharedReg1_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1_out;
SharedReg7_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg7_out;
SharedReg383_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg383_out;
SharedReg290_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg290_out;
SharedReg418_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg418_out;
SharedReg367_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg367_out;
SharedReg480_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg480_out;
   MUX_Subtract4_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg664_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg289_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg290_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg418_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg367_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg480_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg535_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg439_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg367_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg440_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg457_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg7_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg383_out_to_MUX_Subtract4_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract4_2_impl_0_out);

   Delay1No220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_2_impl_0_out,
                 Y => Delay1No220_out);

SharedReg665_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg665_out;
Delay15No17_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_2_cast <= Delay15No17_out;
Delay16No7_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_3_cast <= Delay16No7_out;
SharedReg479_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg479_out;
SharedReg418_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg418_out;
SharedReg418_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg418_out;
SharedReg534_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg534_out;
SharedReg17_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg17_out;
SharedReg23_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg23_out;
SharedReg440_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg440_out;
SharedReg368_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg368_out;
SharedReg479_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg479_out;
SharedReg418_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg418_out;
SharedReg384_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg384_out;
   MUX_Subtract4_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg665_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay15No17_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg368_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg479_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg418_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg384_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => Delay16No7_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg479_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg418_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg418_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg534_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg17_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg23_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg440_out_to_MUX_Subtract4_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract4_2_impl_1_out);

   Delay1No221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_2_impl_1_out,
                 Y => Delay1No221_out);

Delay1No222_out_to_Subtract4_3_impl_parent_implementedSystem_port_0_cast <= Delay1No222_out;
Delay1No223_out_to_Subtract4_3_impl_parent_implementedSystem_port_1_cast <= Delay1No223_out;
   Subtract4_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_3_impl_out,
                 X => Delay1No222_out_to_Subtract4_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No223_out_to_Subtract4_3_impl_parent_implementedSystem_port_1_cast);

SharedReg422_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg422_out;
SharedReg312_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg312_out;
SharedReg484_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg484_out;
SharedReg629_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg629_out;
SharedReg292_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg292_out;
SharedReg539_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg539_out;
SharedReg443_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg443_out;
SharedReg370_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg370_out;
SharedReg444_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg444_out;
SharedReg443_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg443_out;
SharedReg1_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1_out;
SharedReg7_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg7_out;
SharedReg387_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg387_out;
SharedReg293_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg293_out;
   MUX_Subtract4_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg422_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg312_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg7_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg387_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg293_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg484_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg629_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg292_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg539_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg443_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg370_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg444_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg443_out_to_MUX_Subtract4_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract4_3_impl_0_out);

   Delay1No222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_3_impl_0_out,
                 Y => Delay1No222_out);

SharedReg482_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg482_out;
SharedReg403_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg403_out;
SharedReg388_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg388_out;
SharedReg630_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg630_out;
Delay15No18_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_5_cast <= Delay15No18_out;
Delay16No8_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_6_cast <= Delay16No8_out;
SharedReg482_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg482_out;
SharedReg422_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg422_out;
SharedReg422_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg422_out;
SharedReg482_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg482_out;
SharedReg17_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg17_out;
SharedReg23_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg23_out;
SharedReg444_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg444_out;
SharedReg371_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg371_out;
   MUX_Subtract4_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg482_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg403_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg17_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg23_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg444_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg371_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg388_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg630_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay15No18_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay16No8_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg482_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg422_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg422_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg482_out_to_MUX_Subtract4_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract4_3_impl_1_out);

   Delay1No223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_3_impl_1_out,
                 Y => Delay1No223_out);

Delay1No224_out_to_Subtract4_4_impl_parent_implementedSystem_port_0_cast <= Delay1No224_out;
Delay1No225_out_to_Subtract4_4_impl_parent_implementedSystem_port_1_cast <= Delay1No225_out;
   Subtract4_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract4_4_impl_out,
                 X => Delay1No224_out_to_Subtract4_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No225_out_to_Subtract4_4_impl_parent_implementedSystem_port_1_cast);

SharedReg391_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg391_out;
SharedReg322_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg322_out;
SharedReg407_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg407_out;
SharedReg373_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg373_out;
SharedReg448_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg448_out;
SharedReg635_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg635_out;
SharedReg300_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg300_out;
SharedReg543_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg543_out;
SharedReg446_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg446_out;
SharedReg321_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg321_out;
SharedReg427_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg427_out;
SharedReg466_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg466_out;
SharedReg1_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1_out;
SharedReg7_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg7_out;
   MUX_Subtract4_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg391_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg322_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg427_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg466_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg7_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg407_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg373_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg448_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg635_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg300_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg543_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg446_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg321_out_to_MUX_Subtract4_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract4_4_impl_0_out);

   Delay1No224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_4_impl_0_out,
                 Y => Delay1No224_out);

SharedReg447_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg447_out;
SharedReg391_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg391_out;
SharedReg466_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg466_out;
SharedReg426_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg426_out;
SharedReg375_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg375_out;
SharedReg612_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg612_out;
Delay15No19_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_7_cast <= Delay15No19_out;
Delay16No9_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_8_cast <= Delay16No9_out;
SharedReg486_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg486_out;
SharedReg407_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg407_out;
SharedReg426_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg426_out;
SharedReg542_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg542_out;
SharedReg17_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg17_out;
SharedReg23_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg23_out;
   MUX_Subtract4_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg447_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg391_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg426_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg542_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg17_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg23_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg466_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg426_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg375_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg612_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay15No19_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay16No9_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg486_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg407_out_to_MUX_Subtract4_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract4_4_impl_1_out);

   Delay1No225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract4_4_impl_1_out,
                 Y => Delay1No225_out);

Delay1No226_out_to_Product37_0_impl_parent_implementedSystem_port_0_cast <= Delay1No226_out;
Delay1No227_out_to_Product37_0_impl_parent_implementedSystem_port_1_cast <= Delay1No227_out;
   Product37_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product37_0_impl_out,
                 X => Delay1No226_out_to_Product37_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No227_out_to_Product37_0_impl_parent_implementedSystem_port_1_cast);

SharedReg857_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg857_out;
SharedReg835_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg835_out;
SharedReg831_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg831_out;
SharedReg794_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg794_out;
SharedReg36_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg36_out;
SharedReg798_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg798_out;
SharedReg776_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg776_out;
SharedReg705_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg705_out;
SharedReg861_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg861_out;
SharedReg94_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg94_out;
SharedReg736_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg736_out;
SharedReg850_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg850_out;
SharedReg807_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg807_out;
SharedReg833_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg833_out;
   MUX_Product37_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg857_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg835_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg736_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg850_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg807_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg833_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg831_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg794_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg36_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg798_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg776_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg705_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg861_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg94_out_to_MUX_Product37_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product37_0_impl_0_out);

   Delay1No226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_0_impl_0_out,
                 Y => Delay1No226_out);

SharedReg577_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg577_out;
SharedReg704_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg704_out;
SharedReg679_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg679_out;
SharedReg637_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg637_out;
SharedReg819_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg819_out;
SharedReg682_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg682_out;
SharedReg326_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg326_out;
SharedReg853_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg853_out;
SharedReg737_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg737_out;
SharedReg802_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg802_out;
SharedReg826_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg826_out;
SharedReg576_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg576_out;
SharedReg639_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg639_out;
SharedReg704_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg704_out;
   MUX_Product37_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg577_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg704_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg826_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg576_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg639_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg704_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg679_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg637_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg819_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg682_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg326_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg853_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg737_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg802_out_to_MUX_Product37_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product37_0_impl_1_out);

   Delay1No227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_0_impl_1_out,
                 Y => Delay1No227_out);

Delay1No228_out_to_Product37_1_impl_parent_implementedSystem_port_0_cast <= Delay1No228_out;
Delay1No229_out_to_Product37_1_impl_parent_implementedSystem_port_1_cast <= Delay1No229_out;
   Product37_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product37_1_impl_out,
                 X => Delay1No228_out_to_Product37_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No229_out_to_Product37_1_impl_parent_implementedSystem_port_1_cast);

SharedReg850_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg850_out;
SharedReg807_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg807_out;
SharedReg833_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg833_out;
SharedReg857_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg857_out;
SharedReg835_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg835_out;
SharedReg838_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg838_out;
SharedReg794_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg794_out;
SharedReg42_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg42_out;
SharedReg798_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg798_out;
SharedReg776_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg776_out;
SharedReg711_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg711_out;
SharedReg778_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg778_out;
SharedReg779_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg779_out;
SharedReg780_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg780_out;
   MUX_Product37_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg850_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg807_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg711_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg778_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg779_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg780_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg833_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg857_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg835_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg838_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg794_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg42_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg798_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg776_out_to_MUX_Product37_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product37_1_impl_0_out);

   Delay1No228_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_1_impl_0_out,
                 Y => Delay1No228_out);

SharedReg581_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg581_out;
SharedReg644_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg644_out;
SharedReg710_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg710_out;
SharedReg582_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg582_out;
SharedReg710_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg710_out;
SharedReg642_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg642_out;
SharedReg642_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg642_out;
SharedReg819_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg819_out;
SharedReg687_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg687_out;
SharedReg333_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg333_out;
SharedReg853_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg853_out;
SharedReg138_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg138_out;
SharedReg207_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg207_out;
SharedReg115_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg115_out;
   MUX_Product37_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg581_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg644_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg853_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg138_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg207_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg115_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg710_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg582_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg710_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg642_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg642_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg819_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg687_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg333_out_to_MUX_Product37_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product37_1_impl_1_out);

   Delay1No229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_1_impl_1_out,
                 Y => Delay1No229_out);

Delay1No230_out_to_Product37_2_impl_parent_implementedSystem_port_0_cast <= Delay1No230_out;
Delay1No231_out_to_Product37_2_impl_parent_implementedSystem_port_1_cast <= Delay1No231_out;
   Product37_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product37_2_impl_out,
                 X => Delay1No230_out_to_Product37_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No231_out_to_Product37_2_impl_parent_implementedSystem_port_1_cast);

SharedReg861_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg861_out;
SharedReg100_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg100_out;
SharedReg752_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg752_out;
SharedReg824_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg824_out;
SharedReg77_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg77_out;
SharedReg833_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg833_out;
SharedReg852_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg852_out;
SharedReg835_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg835_out;
SharedReg831_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg831_out;
SharedReg74_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg74_out;
SharedReg797_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg797_out;
SharedReg798_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg798_out;
SharedReg776_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg776_out;
SharedReg717_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg717_out;
   MUX_Product37_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg861_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg100_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg797_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg798_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg776_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg717_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg752_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg824_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg77_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg833_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg852_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg835_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg831_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg74_out_to_MUX_Product37_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product37_2_impl_0_out);

   Delay1No230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_2_impl_0_out,
                 Y => Delay1No230_out);

SharedReg753_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg753_out;
SharedReg802_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg802_out;
SharedReg826_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg826_out;
SharedReg753_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg753_out;
SharedReg807_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg807_out;
SharedReg716_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg716_out;
SharedReg587_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg587_out;
SharedReg689_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg689_out;
SharedReg689_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg689_out;
SharedReg816_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg816_out;
SharedReg48_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg48_out;
SharedReg692_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg692_out;
SharedReg340_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg340_out;
SharedReg853_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg853_out;
   MUX_Product37_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg753_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg802_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg48_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg692_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg340_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg853_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg826_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg753_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg807_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg716_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg587_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg689_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg689_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg816_out_to_MUX_Product37_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product37_2_impl_1_out);

   Delay1No231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_2_impl_1_out,
                 Y => Delay1No231_out);

Delay1No232_out_to_Product37_3_impl_parent_implementedSystem_port_0_cast <= Delay1No232_out;
Delay1No233_out_to_Product37_3_impl_parent_implementedSystem_port_1_cast <= Delay1No233_out;
   Product37_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product37_3_impl_out,
                 X => Delay1No232_out_to_Product37_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No233_out_to_Product37_3_impl_parent_implementedSystem_port_1_cast);

SharedReg798_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg798_out;
SharedReg776_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg776_out;
SharedReg723_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg723_out;
SharedReg861_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg861_out;
SharedReg103_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg103_out;
SharedReg780_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg780_out;
SharedReg824_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg824_out;
SharedReg83_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg83_out;
SharedReg833_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg833_out;
SharedReg852_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg852_out;
SharedReg835_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg835_out;
SharedReg838_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg838_out;
SharedReg794_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg794_out;
SharedReg54_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg54_out;
   MUX_Product37_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg798_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg776_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg835_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg838_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg794_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg54_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg723_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg861_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg103_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg780_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg824_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg83_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg833_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg852_out_to_MUX_Product37_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product37_3_impl_0_out);

   Delay1No232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_3_impl_0_out,
                 Y => Delay1No232_out);

SharedReg697_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg697_out;
SharedReg347_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg347_out;
SharedReg853_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg853_out;
SharedReg761_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg761_out;
SharedReg802_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg802_out;
SharedReg125_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg125_out;
SharedReg761_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg761_out;
SharedReg807_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg807_out;
SharedReg722_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg722_out;
SharedReg592_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg592_out;
SharedReg694_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg694_out;
SharedReg652_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg652_out;
SharedReg652_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg652_out;
SharedReg819_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg819_out;
   MUX_Product37_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg697_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg347_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg694_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg652_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg652_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg819_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg853_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg761_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg802_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg125_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg761_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg807_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg722_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg592_out_to_MUX_Product37_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product37_3_impl_1_out);

   Delay1No233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_3_impl_1_out,
                 Y => Delay1No233_out);

Delay1No234_out_to_Product37_4_impl_parent_implementedSystem_port_0_cast <= Delay1No234_out;
Delay1No235_out_to_Product37_4_impl_parent_implementedSystem_port_1_cast <= Delay1No235_out;
   Product37_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product37_4_impl_out,
                 X => Delay1No234_out_to_Product37_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No235_out_to_Product37_4_impl_parent_implementedSystem_port_1_cast);

SharedReg816_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg816_out;
SharedReg60_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg60_out;
SharedReg798_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg798_out;
SharedReg776_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg776_out;
SharedReg729_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg729_out;
SharedReg778_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg778_out;
SharedReg106_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg106_out;
SharedReg768_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg768_out;
SharedReg596_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg596_out;
SharedReg89_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg89_out;
SharedReg127_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg127_out;
SharedReg791_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg791_out;
SharedReg835_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg835_out;
SharedReg831_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg831_out;
   MUX_Product37_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg816_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg60_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg127_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg791_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg835_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg831_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg798_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg776_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg729_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg778_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg106_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg768_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg596_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg89_out_to_MUX_Product37_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product37_4_impl_0_out);

   Delay1No234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_4_impl_0_out,
                 Y => Delay1No234_out);

SharedReg594_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg594_out;
SharedReg819_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg819_out;
SharedReg702_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg702_out;
SharedReg354_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg354_out;
SharedReg853_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg853_out;
SharedReg153_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg153_out;
SharedReg802_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg802_out;
SharedReg826_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg826_out;
SharedReg855_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg855_out;
SharedReg807_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg807_out;
SharedReg813_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg813_out;
SharedReg105_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg105_out;
SharedReg728_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg728_out;
SharedReg699_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg699_out;
   MUX_Product37_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg594_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg819_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg813_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg105_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg728_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg699_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg702_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg354_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg853_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg153_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg802_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg826_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg855_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg807_out_to_MUX_Product37_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product37_4_impl_1_out);

   Delay1No235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product37_4_impl_1_out,
                 Y => Delay1No235_out);

Delay1No236_out_to_Subtract9_0_impl_parent_implementedSystem_port_0_cast <= Delay1No236_out;
Delay1No237_out_to_Subtract9_0_impl_parent_implementedSystem_port_1_cast <= Delay1No237_out;
   Subtract9_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_0_impl_out,
                 X => Delay1No236_out_to_Subtract9_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No237_out_to_Subtract9_0_impl_parent_implementedSystem_port_1_cast);

SharedReg616_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg616_out;
SharedReg2_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg2_out;
SharedReg8_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg8_out;
SharedReg378_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg378_out;
SharedReg672_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg672_out;
SharedReg378_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg378_out;
SharedReg378_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg378_out;
SharedReg410_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg410_out;
SharedReg430_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg430_out;
Delay15No20_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_10_cast <= Delay15No20_out;
SharedReg245_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg245_out;
SharedReg671_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg671_out;
SharedReg470_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg470_out;
SharedReg430_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg430_out;
   MUX_Subtract9_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg616_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg2_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg245_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg671_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg470_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg430_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg8_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg378_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg672_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg378_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg378_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg410_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg430_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay15No20_out_to_MUX_Subtract9_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract9_0_impl_0_out);

   Delay1No236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_0_impl_0_out,
                 Y => Delay1No236_out);

SharedReg634_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg634_out;
SharedReg18_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg18_out;
SharedReg24_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg24_out;
SharedReg432_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg432_out;
SharedReg620_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg620_out;
SharedReg671_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg671_out;
SharedReg453_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg453_out;
SharedReg470_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg470_out;
SharedReg394_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg394_out;
SharedReg526_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg526_out;
SharedReg204_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg204_out;
SharedReg286_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg286_out;
SharedReg378_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg378_out;
SharedReg525_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg525_out;
   MUX_Subtract9_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg634_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg18_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg204_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg286_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg378_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg525_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg24_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg432_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg620_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg671_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg453_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg470_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg394_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg526_out_to_MUX_Subtract9_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract9_0_impl_1_out);

   Delay1No237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_0_impl_1_out,
                 Y => Delay1No237_out);

Delay1No238_out_to_Subtract9_1_impl_parent_implementedSystem_port_0_cast <= Delay1No238_out;
Delay1No239_out_to_Subtract9_1_impl_parent_implementedSystem_port_1_cast <= Delay1No239_out;
   Subtract9_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_1_impl_out,
                 X => Delay1No238_out_to_Subtract9_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No239_out_to_Subtract9_1_impl_parent_implementedSystem_port_1_cast);

SharedReg674_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg674_out;
SharedReg454_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg454_out;
SharedReg414_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg414_out;
SharedReg529_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg529_out;
SharedReg2_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg2_out;
SharedReg8_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg8_out;
SharedReg381_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg381_out;
SharedReg675_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg675_out;
SharedReg381_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg381_out;
SharedReg381_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg381_out;
SharedReg414_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg414_out;
SharedReg435_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg435_out;
Delay15No21_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_13_cast <= Delay15No21_out;
SharedReg254_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg254_out;
   MUX_Subtract9_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg674_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg454_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg414_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg435_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay15No21_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg254_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg414_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg529_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg2_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg8_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg381_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg675_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg381_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg381_out_to_MUX_Subtract9_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract9_1_impl_0_out);

   Delay1No238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_1_impl_0_out,
                 Y => Delay1No238_out);

SharedReg289_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg289_out;
SharedReg381_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg381_out;
SharedReg475_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg475_out;
SharedReg623_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg623_out;
SharedReg18_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg18_out;
SharedReg24_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg24_out;
SharedReg437_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg437_out;
SharedReg625_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg625_out;
SharedReg674_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg674_out;
SharedReg456_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg456_out;
SharedReg475_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg475_out;
SharedReg397_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg397_out;
SharedReg530_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg530_out;
SharedReg212_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg212_out;
   MUX_Subtract9_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg289_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg381_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg475_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg397_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg530_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg212_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg475_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg623_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg18_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg24_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg437_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg625_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg674_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg456_out_to_MUX_Subtract9_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract9_1_impl_1_out);

   Delay1No239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_1_impl_1_out,
                 Y => Delay1No239_out);

Delay1No240_out_to_Subtract9_2_impl_parent_implementedSystem_port_0_cast <= Delay1No240_out;
Delay1No241_out_to_Subtract9_2_impl_parent_implementedSystem_port_1_cast <= Delay1No241_out;
   Subtract9_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_2_impl_out,
                 X => Delay1No240_out_to_Subtract9_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No241_out_to_Subtract9_2_impl_parent_implementedSystem_port_1_cast);

SharedReg457_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg457_out;
Delay15No22_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_2_cast <= Delay15No22_out;
SharedReg263_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg263_out;
SharedReg665_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg665_out;
SharedReg479_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg479_out;
SharedReg439_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg439_out;
SharedReg599_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg599_out;
SharedReg2_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg2_out;
SharedReg8_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg8_out;
SharedReg402_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg402_out;
SharedReg573_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg573_out;
SharedReg384_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg384_out;
SharedReg402_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg402_out;
SharedReg439_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg439_out;
   MUX_Subtract9_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg457_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay15No22_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg573_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg384_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg402_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg439_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg263_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg665_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg479_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg439_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg599_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg2_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg8_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg402_out_to_MUX_Subtract9_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract9_2_impl_0_out);

   Delay1No240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_2_impl_0_out,
                 Y => Delay1No240_out);

SharedReg419_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg419_out;
SharedReg600_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg600_out;
SharedReg220_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg220_out;
SharedReg571_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg571_out;
SharedReg384_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg384_out;
SharedReg534_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg534_out;
SharedReg628_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg628_out;
SharedReg18_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg18_out;
SharedReg24_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg24_out;
SharedReg459_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg459_out;
SharedReg604_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg604_out;
SharedReg572_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg572_out;
SharedReg481_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg481_out;
SharedReg534_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg534_out;
   MUX_Subtract9_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg419_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg600_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg604_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg572_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg481_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg534_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg220_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg571_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg384_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg534_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg628_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg18_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg24_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg459_out_to_MUX_Subtract9_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract9_2_impl_1_out);

   Delay1No241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_2_impl_1_out,
                 Y => Delay1No241_out);

Delay1No242_out_to_Subtract9_3_impl_parent_implementedSystem_port_0_cast <= Delay1No242_out;
Delay1No243_out_to_Subtract9_3_impl_parent_implementedSystem_port_1_cast <= Delay1No243_out;
   Subtract9_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_3_impl_out,
                 X => Delay1No242_out_to_Subtract9_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No243_out_to_Subtract9_3_impl_parent_implementedSystem_port_1_cast);

SharedReg388_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg388_out;
SharedReg405_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg405_out;
SharedReg422_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg422_out;
SharedReg443_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg443_out;
Delay15No23_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_5_cast <= Delay15No23_out;
SharedReg272_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg272_out;
SharedReg668_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg668_out;
SharedReg482_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg482_out;
SharedReg443_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg443_out;
SharedReg538_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg538_out;
SharedReg2_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg2_out;
SharedReg8_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg8_out;
SharedReg405_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg405_out;
SharedReg296_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg296_out;
   MUX_Subtract9_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg388_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg405_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg2_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg8_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg405_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg296_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg422_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg443_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay15No23_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg272_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg668_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg482_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg443_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg538_out_to_MUX_Subtract9_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract9_3_impl_0_out);

   Delay1No242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_3_impl_0_out,
                 Y => Delay1No242_out);

SharedReg295_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg295_out;
SharedReg485_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg485_out;
SharedReg482_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg482_out;
SharedReg404_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg404_out;
SharedReg539_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg539_out;
SharedReg228_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg228_out;
SharedReg294_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg294_out;
SharedReg388_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg388_out;
SharedReg538_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg538_out;
SharedReg631_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg631_out;
SharedReg18_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg18_out;
SharedReg24_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg24_out;
SharedReg463_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg463_out;
SharedReg610_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg610_out;
   MUX_Subtract9_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg295_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg485_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg18_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg24_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg463_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg610_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg482_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg404_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg539_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg228_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg294_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg388_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg538_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg631_out_to_MUX_Subtract9_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract9_3_impl_1_out);

   Delay1No243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_3_impl_1_out,
                 Y => Delay1No243_out);

Delay1No244_out_to_Subtract9_4_impl_parent_implementedSystem_port_0_cast <= Delay1No244_out;
Delay1No245_out_to_Subtract9_4_impl_parent_implementedSystem_port_1_cast <= Delay1No245_out;
   Subtract9_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract9_4_impl_out,
                 X => Delay1No244_out_to_Subtract9_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No245_out_to_Subtract9_4_impl_parent_implementedSystem_port_1_cast);

SharedReg375_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg375_out;
Delay3No249_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_2_cast <= Delay3No249_out;
SharedReg409_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg409_out;
SharedReg375_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg375_out;
SharedReg407_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg407_out;
SharedReg446_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg446_out;
Delay15No24_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_7_cast <= Delay15No24_out;
SharedReg281_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg281_out;
SharedReg677_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg677_out;
SharedReg466_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg466_out;
SharedReg446_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg446_out;
SharedReg611_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg611_out;
SharedReg2_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg2_out;
SharedReg8_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg8_out;
   MUX_Subtract9_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg375_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay3No249_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg446_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg611_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg2_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg8_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg409_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg375_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg407_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg446_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay15No24_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg281_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg677_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg466_out_to_MUX_Subtract9_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract9_4_impl_0_out);

   Delay1No244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_4_impl_0_out,
                 Y => Delay1No244_out);

SharedReg428_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg428_out;
SharedReg615_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg615_out;
SharedReg636_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg636_out;
SharedReg489_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg489_out;
SharedReg466_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg466_out;
SharedReg391_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg391_out;
SharedReg543_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg543_out;
SharedReg236_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg236_out;
SharedReg734_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg734_out;
SharedReg392_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg392_out;
SharedReg542_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg542_out;
SharedReg613_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg613_out;
SharedReg18_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg18_out;
SharedReg24_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg24_out;
   MUX_Subtract9_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg428_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg615_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg542_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg613_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg18_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg24_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg636_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg489_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg466_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg391_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg543_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg236_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg734_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg392_out_to_MUX_Subtract9_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract9_4_impl_1_out);

   Delay1No245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract9_4_impl_1_out,
                 Y => Delay1No245_out);

Delay1No246_out_to_Product39_3_impl_parent_implementedSystem_port_0_cast <= Delay1No246_out;
Delay1No247_out_to_Product39_3_impl_parent_implementedSystem_port_1_cast <= Delay1No247_out;
   Product39_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product39_3_impl_out,
                 X => Delay1No246_out_to_Product39_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No247_out_to_Product39_3_impl_parent_implementedSystem_port_1_cast);

SharedReg257_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg257_out;
SharedReg779_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg779_out;
SharedReg803_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg803_out;
SharedReg855_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg855_out;
SharedReg781_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg781_out;
SharedReg80_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg80_out;
SharedReg690_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg690_out;
SharedReg835_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg835_out;
SharedReg843_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg843_out;
SharedReg794_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg794_out;
SharedReg795_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg795_out;
SharedReg787_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg787_out;
SharedReg862_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg862_out;
SharedReg585_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg585_out;
   MUX_Product39_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg257_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg779_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg795_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg787_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg862_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg585_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg803_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg855_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg781_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg80_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg690_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg835_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg843_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg794_out_to_MUX_Product39_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product39_3_impl_0_out);

   Delay1No246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product39_3_impl_0_out,
                 Y => Delay1No246_out);

SharedReg801_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg801_out;
SharedReg258_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg258_out;
SharedReg175_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg175_out;
SharedReg718_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg718_out;
SharedReg47_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg47_out;
SharedReg805_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg805_out;
SharedReg841_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg841_out;
SharedReg647_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg647_out;
SharedReg716_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg716_out;
SharedReg689_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg689_out;
SharedReg754_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg754_out;
Delay9No3_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_12_cast <= Delay9No3_out;
SharedReg584_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg584_out;
SharedReg863_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg863_out;
   MUX_Product39_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg801_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg258_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg754_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay9No3_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg584_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg863_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg175_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg718_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg47_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg805_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg841_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg647_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg716_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg689_out_to_MUX_Product39_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product39_3_impl_1_out);

   Delay1No247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product39_3_impl_1_out,
                 Y => Delay1No247_out);

Delay1No248_out_to_Subtract20_0_impl_parent_implementedSystem_port_0_cast <= Delay1No248_out;
Delay1No249_out_to_Subtract20_0_impl_parent_implementedSystem_port_1_cast <= Delay1No249_out;
   Subtract20_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract20_0_impl_out,
                 X => Delay1No248_out_to_Subtract20_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No249_out_to_Subtract20_0_impl_parent_implementedSystem_port_1_cast);

SharedReg670_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg670_out;
SharedReg3_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg3_out;
SharedReg9_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg9_out;
SharedReg634_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg634_out;
SharedReg197_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg197_out;
SharedReg547_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg547_out;
SharedReg412_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg412_out;
SharedReg550_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg550_out;
SharedReg670_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg670_out;
Delay15No30_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_10_cast <= Delay15No30_out;
SharedReg525_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg525_out;
SharedReg203_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg203_out;
SharedReg326_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg326_out;
SharedReg670_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg670_out;
   MUX_Subtract20_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg670_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg3_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg525_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg203_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg326_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg670_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg9_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg634_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg197_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg547_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg412_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg550_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg670_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay15No30_out_to_MUX_Subtract20_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract20_0_impl_0_out);

   Delay1No248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_0_impl_0_out,
                 Y => Delay1No248_out);

SharedReg633_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg633_out;
SharedReg19_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg19_out;
SharedReg25_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg25_out;
SharedReg633_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg633_out;
SharedReg237_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg237_out;
SharedReg575_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg575_out;
SharedReg474_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg474_out;
SharedReg496_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg496_out;
SharedReg287_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg287_out;
SharedReg470_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg470_out;
SharedReg632_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg632_out;
SharedReg237_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg237_out;
SharedReg491_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg491_out;
SharedReg287_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg287_out;
   MUX_Subtract20_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg633_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg19_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg632_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg237_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg491_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg287_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg25_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg633_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg237_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg575_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg474_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg496_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg287_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg470_out_to_MUX_Subtract20_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract20_0_impl_1_out);

   Delay1No249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_0_impl_1_out,
                 Y => Delay1No249_out);

Delay1No250_out_to_Subtract20_1_impl_parent_implementedSystem_port_0_cast <= Delay1No250_out;
Delay1No251_out_to_Subtract20_1_impl_parent_implementedSystem_port_1_cast <= Delay1No251_out;
   Subtract20_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract20_1_impl_out,
                 X => Delay1No250_out_to_Subtract20_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No251_out_to_Subtract20_1_impl_parent_implementedSystem_port_1_cast);

SharedReg211_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg211_out;
SharedReg333_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg333_out;
SharedReg662_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg662_out;
SharedReg662_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg662_out;
SharedReg3_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg3_out;
SharedReg9_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg9_out;
Delay3No206_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_7_cast <= Delay3No206_out;
SharedReg205_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg205_out;
SharedReg552_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg552_out;
SharedReg416_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg416_out;
SharedReg555_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg555_out;
SharedReg673_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg673_out;
Delay15No31_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_13_cast <= Delay15No31_out;
SharedReg529_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg529_out;
   MUX_Subtract20_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg211_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg333_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg555_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg673_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay15No31_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg529_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg662_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg662_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg3_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg9_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay3No206_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg205_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg552_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg416_out_to_MUX_Subtract20_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract20_1_impl_0_out);

   Delay1No250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_1_impl_0_out,
                 Y => Delay1No250_out);

SharedReg246_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg246_out;
SharedReg498_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg498_out;
SharedReg674_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg674_out;
SharedReg622_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg622_out;
SharedReg19_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg19_out;
SharedReg25_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg25_out;
SharedReg663_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg663_out;
SharedReg246_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg246_out;
SharedReg580_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg580_out;
SharedReg478_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg478_out;
SharedReg503_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg503_out;
SharedReg290_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg290_out;
SharedReg475_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg475_out;
SharedReg662_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg662_out;
   MUX_Subtract20_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg246_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg498_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg503_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg290_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg475_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg662_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg674_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg622_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg19_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg25_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg663_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg246_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg580_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg478_out_to_MUX_Subtract20_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract20_1_impl_1_out);

   Delay1No251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_1_impl_1_out,
                 Y => Delay1No251_out);

Delay1No252_out_to_Subtract20_2_impl_parent_implementedSystem_port_0_cast <= Delay1No252_out;
Delay1No253_out_to_Subtract20_2_impl_parent_implementedSystem_port_1_cast <= Delay1No253_out;
   Subtract20_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract20_2_impl_out,
                 X => Delay1No252_out_to_Subtract20_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No253_out_to_Subtract20_2_impl_parent_implementedSystem_port_1_cast);

SharedReg571_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg571_out;
Delay15No32_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_2_cast <= Delay15No32_out;
SharedReg534_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg534_out;
SharedReg219_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg219_out;
SharedReg340_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg340_out;
SharedReg664_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg664_out;
SharedReg664_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg664_out;
SharedReg3_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg3_out;
SharedReg9_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg9_out;
SharedReg666_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg666_out;
SharedReg213_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg213_out;
SharedReg557_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg557_out;
SharedReg441_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg441_out;
SharedReg560_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg560_out;
   MUX_Subtract20_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg571_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay15No32_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg213_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg557_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg441_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg560_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg534_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg219_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg340_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg664_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg664_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg3_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg9_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg666_out_to_MUX_Subtract20_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract20_2_impl_0_out);

   Delay1No252_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_2_impl_0_out,
                 Y => Delay1No252_out);

SharedReg293_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg293_out;
SharedReg479_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg479_out;
SharedReg626_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg626_out;
SharedReg255_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg255_out;
SharedReg505_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg505_out;
SharedReg572_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg572_out;
SharedReg627_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg627_out;
SharedReg19_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg19_out;
SharedReg25_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg25_out;
SharedReg665_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg665_out;
SharedReg255_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg255_out;
SharedReg585_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg585_out;
SharedReg537_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg537_out;
SharedReg510_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg510_out;
   MUX_Subtract20_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg293_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg479_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg255_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg585_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg537_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg510_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg626_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg255_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg505_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg572_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg627_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg19_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg25_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg665_out_to_MUX_Subtract20_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract20_2_impl_1_out);

   Delay1No253_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_2_impl_1_out,
                 Y => Delay1No253_out);

Delay1No254_out_to_Subtract20_3_impl_parent_implementedSystem_port_0_cast <= Delay1No254_out;
Delay1No255_out_to_Subtract20_3_impl_parent_implementedSystem_port_1_cast <= Delay1No255_out;
   Subtract20_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract20_3_impl_out,
                 X => Delay1No254_out_to_Subtract20_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No255_out_to_Subtract20_3_impl_parent_implementedSystem_port_1_cast);

SharedReg562_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg562_out;
SharedReg445_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg445_out;
SharedReg565_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg565_out;
SharedReg667_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg667_out;
Delay15No33_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_5_cast <= Delay15No33_out;
SharedReg538_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg538_out;
SharedReg227_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg227_out;
SharedReg347_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg347_out;
SharedReg667_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg667_out;
SharedReg629_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg629_out;
SharedReg3_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg3_out;
SharedReg9_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg9_out;
SharedReg669_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg669_out;
SharedReg221_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg221_out;
   MUX_Subtract20_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg562_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg445_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg3_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg9_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg669_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg221_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg565_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg667_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay15No33_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg538_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg227_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg347_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg667_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg629_out_to_MUX_Subtract20_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract20_3_impl_0_out);

   Delay1No254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_3_impl_0_out,
                 Y => Delay1No254_out);

SharedReg590_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg590_out;
SharedReg541_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg541_out;
SharedReg517_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg517_out;
SharedReg295_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg295_out;
SharedReg482_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg482_out;
SharedReg629_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg629_out;
SharedReg264_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg264_out;
SharedReg512_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg512_out;
SharedReg295_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg295_out;
SharedReg630_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg630_out;
SharedReg19_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg19_out;
SharedReg25_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg25_out;
SharedReg668_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg668_out;
SharedReg264_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg264_out;
   MUX_Subtract20_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg590_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg541_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg19_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg25_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg668_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg264_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg517_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg295_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg482_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg629_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg264_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg512_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg295_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg630_out_to_MUX_Subtract20_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract20_3_impl_1_out);

   Delay1No255_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_3_impl_1_out,
                 Y => Delay1No255_out);

Delay1No256_out_to_Subtract20_4_impl_parent_implementedSystem_port_0_cast <= Delay1No256_out;
Delay1No257_out_to_Subtract20_4_impl_parent_implementedSystem_port_1_cast <= Delay1No257_out;
   Subtract20_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract20_4_impl_out,
                 X => Delay1No256_out_to_Subtract20_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No257_out_to_Subtract20_4_impl_parent_implementedSystem_port_1_cast);

SharedReg613_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg613_out;
SharedReg229_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg229_out;
SharedReg567_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg567_out;
SharedReg409_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg409_out;
SharedReg570_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg570_out;
SharedReg676_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg676_out;
Delay15No34_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_7_cast <= Delay15No34_out;
SharedReg542_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg542_out;
SharedReg235_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg235_out;
SharedReg354_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg354_out;
SharedReg676_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg676_out;
SharedReg676_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg676_out;
SharedReg3_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg3_out;
SharedReg9_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg9_out;
   MUX_Subtract20_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg613_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg229_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg676_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg676_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg3_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg9_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg567_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg409_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg570_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg676_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay15No34_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg542_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg235_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg354_out_to_MUX_Subtract20_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract20_4_impl_0_out);

   Delay1No256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_4_impl_0_out,
                 Y => Delay1No256_out);

SharedReg677_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg677_out;
SharedReg273_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg273_out;
SharedReg595_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg595_out;
SharedReg545_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg545_out;
SharedReg524_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg524_out;
SharedReg677_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg677_out;
SharedReg486_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg486_out;
SharedReg635_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg635_out;
SharedReg273_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg273_out;
SharedReg519_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg519_out;
SharedReg677_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg677_out;
SharedReg636_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg636_out;
SharedReg19_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg19_out;
SharedReg25_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg25_out;
   MUX_Subtract20_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg677_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg273_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg677_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg636_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg19_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg25_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg595_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg545_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg524_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg677_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg486_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg635_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg273_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg519_out_to_MUX_Subtract20_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract20_4_impl_1_out);

   Delay1No257_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract20_4_impl_1_out,
                 Y => Delay1No257_out);

Delay1No258_out_to_Product220_2_impl_parent_implementedSystem_port_0_cast <= Delay1No258_out;
Delay1No259_out_to_Product220_2_impl_parent_implementedSystem_port_1_cast <= Delay1No259_out;
   Product220_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product220_2_impl_out,
                 X => Delay1No258_out_to_Product220_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No259_out_to_Product220_2_impl_parent_implementedSystem_port_1_cast);

SharedReg778_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg778_out;
SharedReg779_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg779_out;
SharedReg780_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg780_out;
SharedReg850_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg850_out;
SharedReg807_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg807_out;
SharedReg833_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg833_out;
SharedReg857_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg857_out;
SharedReg835_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg835_out;
SharedReg838_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg838_out;
SharedReg794_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg794_out;
SharedReg48_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg48_out;
SharedReg796_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg796_out;
SharedReg799_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg799_out;
SharedReg214_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg214_out;
   MUX_Product220_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg778_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg779_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg48_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg796_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg799_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg214_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg780_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg850_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg807_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg833_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg857_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg835_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg838_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg794_out_to_MUX_Product220_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product220_2_impl_0_out);

   Delay1No258_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product220_2_impl_0_out,
                 Y => Delay1No258_out);

SharedReg143_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg143_out;
SharedReg215_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg215_out;
SharedReg120_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg120_out;
SharedReg586_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg586_out;
SharedReg649_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg649_out;
SharedReg752_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg752_out;
SharedReg587_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg587_out;
SharedReg716_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg716_out;
SharedReg647_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg647_out;
SharedReg647_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg647_out;
SharedReg819_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg819_out;
SharedReg647_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg647_out;
SharedReg340_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg340_out;
SharedReg800_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg800_out;
   MUX_Product220_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg143_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg215_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg819_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg647_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg340_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg800_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg120_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg586_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg649_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg752_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg587_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg716_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg647_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg647_out_to_MUX_Product220_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product220_2_impl_1_out);

   Delay1No259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product220_2_impl_1_out,
                 Y => Delay1No259_out);

Delay1No260_out_to_Product220_3_impl_parent_implementedSystem_port_0_cast <= Delay1No260_out;
Delay1No261_out_to_Product220_3_impl_parent_implementedSystem_port_1_cast <= Delay1No261_out;
   Product220_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product220_3_impl_out,
                 X => Delay1No260_out_to_Product220_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No261_out_to_Product220_3_impl_parent_implementedSystem_port_1_cast);

SharedReg796_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg796_out;
SharedReg799_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg799_out;
SharedReg222_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg222_out;
SharedReg778_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg778_out;
SharedReg779_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg779_out;
SharedReg803_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg803_out;
SharedReg850_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg850_out;
SharedReg807_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg807_out;
SharedReg833_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg833_out;
SharedReg857_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg857_out;
SharedReg835_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg835_out;
SharedReg694_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg694_out;
SharedReg816_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg816_out;
SharedReg797_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg797_out;
   MUX_Product220_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg796_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg799_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg835_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg694_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg816_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg797_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg222_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg778_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg779_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg803_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg850_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg807_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg833_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg857_out_to_MUX_Product220_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product220_3_impl_0_out);

   Delay1No260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product220_3_impl_0_out,
                 Y => Delay1No260_out);

SharedReg652_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg652_out;
SharedReg347_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg347_out;
SharedReg800_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg800_out;
SharedReg148_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg148_out;
SharedReg223_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg223_out;
SharedReg125_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg125_out;
SharedReg591_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg591_out;
SharedReg654_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg654_out;
SharedReg760_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg760_out;
SharedReg592_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg592_out;
SharedReg722_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg722_out;
SharedReg838_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg838_out;
SharedReg589_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg589_out;
SharedReg765_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg765_out;
   MUX_Product220_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg652_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg347_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg722_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg838_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg589_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg765_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg800_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg148_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg223_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg125_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg591_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg654_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg760_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg592_out_to_MUX_Product220_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product220_3_impl_1_out);

   Delay1No261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product220_3_impl_1_out,
                 Y => Delay1No261_out);

Delay1No262_out_to_Product220_4_impl_parent_implementedSystem_port_0_cast <= Delay1No262_out;
Delay1No263_out_to_Product220_4_impl_parent_implementedSystem_port_1_cast <= Delay1No263_out;
   Product220_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product220_4_impl_out,
                 X => Delay1No262_out_to_Product220_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No263_out_to_Product220_4_impl_parent_implementedSystem_port_1_cast);

SharedReg657_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg657_out;
SharedReg797_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg797_out;
SharedReg796_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg796_out;
SharedReg799_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg799_out;
SharedReg230_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg230_out;
SharedReg153_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg153_out;
SharedReg779_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg779_out;
SharedReg780_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg780_out;
SharedReg850_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg850_out;
SharedReg807_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg807_out;
SharedReg833_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg833_out;
SharedReg834_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg834_out;
SharedReg842_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg842_out;
SharedReg838_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg838_out;
   MUX_Product220_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg657_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg797_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg833_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg834_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg842_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg838_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg796_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg799_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg230_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg153_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg779_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg780_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg850_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg807_out_to_MUX_Product220_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product220_4_impl_0_out);

   Delay1No262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product220_4_impl_0_out,
                 Y => Delay1No262_out);

SharedReg816_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg816_out;
SharedReg773_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg773_out;
SharedReg657_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg657_out;
SharedReg354_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg354_out;
SharedReg800_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg800_out;
SharedReg801_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg801_out;
SharedReg231_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg231_out;
SharedReg130_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg130_out;
SharedReg730_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg730_out;
SharedReg659_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg659_out;
SharedReg728_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg728_out;
SharedReg700_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg700_out;
SharedReg699_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg699_out;
SharedReg657_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg657_out;
   MUX_Product220_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg816_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg773_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg728_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg700_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg699_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg657_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg657_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg354_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg800_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg801_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg231_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg130_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg730_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg659_out_to_MUX_Product220_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product220_4_impl_1_out);

   Delay1No263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product220_4_impl_1_out,
                 Y => Delay1No263_out);

Delay1No264_out_to_Product323_0_impl_parent_implementedSystem_port_0_cast <= Delay1No264_out;
Delay1No265_out_to_Product323_0_impl_parent_implementedSystem_port_1_cast <= Delay1No265_out;
   Product323_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product323_0_impl_out,
                 X => Delay1No264_out_to_Product323_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No265_out_to_Product323_0_impl_parent_implementedSystem_port_1_cast);

SharedReg791_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg791_out;
SharedReg842_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg842_out;
SharedReg838_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg838_out;
SharedReg816_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg816_out;
SharedReg797_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg797_out;
SharedReg796_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg796_out;
SharedReg799_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg799_out;
SharedReg198_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg198_out;
SharedReg778_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg778_out;
SharedReg779_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg779_out;
SharedReg780_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg780_out;
SharedReg576_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg576_out;
SharedReg851_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg851_out;
SharedReg833_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg833_out;
   MUX_Product323_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg791_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg842_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg780_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg576_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg851_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg833_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg838_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg816_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg797_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg796_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg799_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg198_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg778_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg779_out_to_MUX_Product323_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product323_0_impl_0_out);

   Delay1No264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_0_impl_0_out,
                 Y => Delay1No264_out);

SharedReg93_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg93_out;
SharedReg679_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg679_out;
SharedReg637_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg637_out;
SharedReg574_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg574_out;
SharedReg741_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg741_out;
SharedReg637_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg637_out;
SharedReg326_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg326_out;
SharedReg800_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg800_out;
SharedReg133_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg133_out;
SharedReg199_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg199_out;
SharedReg110_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg110_out;
SharedReg855_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg855_out;
SharedReg739_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg739_out;
SharedReg736_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg736_out;
   MUX_Product323_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg93_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg679_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg110_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg855_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg739_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg736_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg637_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg574_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg741_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg637_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg326_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg800_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg133_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg199_out_to_MUX_Product323_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product323_0_impl_1_out);

   Delay1No265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_0_impl_1_out,
                 Y => Delay1No265_out);

Delay1No266_out_to_Product323_1_impl_parent_implementedSystem_port_0_cast <= Delay1No266_out;
Delay1No267_out_to_Product323_1_impl_parent_implementedSystem_port_1_cast <= Delay1No267_out;
   Product323_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product323_1_impl_out,
                 X => Delay1No266_out_to_Product323_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No267_out_to_Product323_1_impl_parent_implementedSystem_port_1_cast);

SharedReg581_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg581_out;
SharedReg851_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg851_out;
SharedReg833_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg833_out;
SharedReg791_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg791_out;
SharedReg842_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg842_out;
SharedReg684_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg684_out;
SharedReg816_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg816_out;
SharedReg797_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg797_out;
SharedReg796_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg796_out;
SharedReg799_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg799_out;
SharedReg206_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg206_out;
SharedReg138_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg138_out;
SharedReg207_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg207_out;
SharedReg803_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg803_out;
   MUX_Product323_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg581_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg851_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg206_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg138_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg207_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg803_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg833_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg791_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg842_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg684_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg816_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg797_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg796_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg799_out_to_MUX_Product323_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product323_1_impl_0_out);

   Delay1No266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_1_impl_0_out,
                 Y => Delay1No266_out);

SharedReg855_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg855_out;
SharedReg747_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg747_out;
SharedReg744_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg744_out;
SharedReg96_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg96_out;
SharedReg684_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg684_out;
SharedReg838_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg838_out;
SharedReg579_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg579_out;
SharedReg749_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg749_out;
SharedReg642_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg642_out;
SharedReg333_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg333_out;
SharedReg800_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg800_out;
SharedReg801_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg801_out;
SharedReg802_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg802_out;
SharedReg115_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg115_out;
   MUX_Product323_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg855_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg747_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg800_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg801_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg802_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg115_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg744_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg96_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg684_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg838_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg579_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg749_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg642_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg333_out_to_MUX_Product323_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product323_1_impl_1_out);

   Delay1No267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_1_impl_1_out,
                 Y => Delay1No267_out);

Delay1No268_out_to_Product323_2_impl_parent_implementedSystem_port_0_cast <= Delay1No268_out;
Delay1No269_out_to_Product323_2_impl_parent_implementedSystem_port_1_cast <= Delay1No269_out;
   Product323_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product323_2_impl_out,
                 X => Delay1No268_out_to_Product323_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No269_out_to_Product323_2_impl_parent_implementedSystem_port_1_cast);

SharedReg143_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg143_out;
SharedReg215_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg215_out;
SharedReg803_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg803_out;
SharedReg586_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg586_out;
SharedReg851_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg851_out;
SharedReg840_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg840_out;
SharedReg791_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg791_out;
SharedReg842_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg842_out;
SharedReg689_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg689_out;
SharedReg816_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg816_out;
SharedReg797_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg797_out;
SharedReg820_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg820_out;
SharedReg504_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg504_out;
SharedReg777_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg777_out;
   MUX_Product323_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg143_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg215_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg797_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg820_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg504_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg777_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg803_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg586_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg851_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg840_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg791_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg842_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg689_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg816_out_to_MUX_Product323_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product323_2_impl_0_out);

   Delay1No268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_2_impl_0_out,
                 Y => Delay1No268_out);

SharedReg801_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg801_out;
SharedReg802_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg802_out;
SharedReg120_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg120_out;
SharedReg855_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg855_out;
SharedReg755_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg755_out;
SharedReg716_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg716_out;
SharedReg99_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg99_out;
SharedReg689_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg689_out;
SharedReg838_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg838_out;
SharedReg584_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg584_out;
SharedReg757_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg757_out;
SharedReg692_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg692_out;
SharedReg799_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg799_out;
SharedReg505_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg505_out;
   MUX_Product323_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg801_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg802_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg757_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg692_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg799_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg505_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg120_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg855_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg755_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg716_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg99_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg689_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg838_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg584_out_to_MUX_Product323_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product323_2_impl_1_out);

   Delay1No269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_2_impl_1_out,
                 Y => Delay1No269_out);

Delay1No270_out_to_Product323_3_impl_parent_implementedSystem_port_0_cast <= Delay1No270_out;
Delay1No271_out_to_Product323_3_impl_parent_implementedSystem_port_1_cast <= Delay1No271_out;
   Product323_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product323_3_impl_out,
                 X => Delay1No270_out_to_Product323_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No271_out_to_Product323_3_impl_parent_implementedSystem_port_1_cast);

SharedReg820_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg820_out;
SharedReg511_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg511_out;
SharedReg777_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg777_out;
SharedReg148_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg148_out;
SharedReg223_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg223_out;
SharedReg780_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg780_out;
SharedReg591_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg591_out;
SharedReg851_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg851_out;
SharedReg840_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg840_out;
SharedReg791_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg791_out;
SharedReg842_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg842_out;
SharedReg836_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg836_out;
SharedReg652_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg652_out;
SharedReg795_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg795_out;
   MUX_Product323_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg820_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg511_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg842_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg836_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg652_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg795_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg777_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg148_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg223_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg780_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg591_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg851_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg840_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg791_out_to_MUX_Product323_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product323_3_impl_0_out);

   Delay1No270_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_3_impl_0_out,
                 Y => Delay1No270_out);

SharedReg697_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg697_out;
SharedReg799_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg799_out;
SharedReg512_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg512_out;
SharedReg801_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg801_out;
SharedReg802_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg802_out;
SharedReg183_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg183_out;
SharedReg855_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg855_out;
SharedReg763_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg763_out;
SharedReg722_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg722_out;
SharedReg102_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg102_out;
SharedReg694_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg694_out;
SharedReg722_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg722_out;
SharedReg816_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg816_out;
SharedReg590_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg590_out;
   MUX_Product323_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg697_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg799_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg694_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg722_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg816_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg590_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg512_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg801_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg802_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg183_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg855_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg763_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg722_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg102_out_to_MUX_Product323_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product323_3_impl_1_out);

   Delay1No271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product323_3_impl_1_out,
                 Y => Delay1No271_out);

Delay1No272_out_to_Product325_0_impl_parent_implementedSystem_port_0_cast <= Delay1No272_out;
Delay1No273_out_to_Product325_0_impl_parent_implementedSystem_port_1_cast <= Delay1No273_out;
   Product325_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product325_0_impl_out,
                 X => Delay1No272_out_to_Product325_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No273_out_to_Product325_0_impl_parent_implementedSystem_port_1_cast);

SharedReg834_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg834_out;
SharedReg704_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg704_out;
SharedReg679_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg679_out;
SharedReg637_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg637_out;
SharedReg795_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg795_out;
SharedReg820_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg820_out;
SharedReg490_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg490_out;
SharedReg777_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg777_out;
SharedReg133_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg133_out;
SharedReg199_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg199_out;
SharedReg803_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg803_out;
SharedReg850_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg850_out;
SharedReg739_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg739_out;
SharedReg840_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg840_out;
   MUX_Product325_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg834_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg704_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg803_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg850_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg739_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg840_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg679_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg637_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg795_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg820_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg490_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg777_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg133_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg199_out_to_MUX_Product325_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product325_0_impl_0_out);

   Delay1No272_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product325_0_impl_0_out,
                 Y => Delay1No272_out);

SharedReg680_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg680_out;
SharedReg842_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg842_out;
SharedReg838_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg838_out;
SharedReg816_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg816_out;
SharedReg575_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg575_out;
SharedReg682_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg682_out;
SharedReg799_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg799_out;
SharedReg491_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg491_out;
SharedReg801_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg801_out;
SharedReg802_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg802_out;
SharedReg110_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg110_out;
SharedReg706_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg706_out;
SharedReg856_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg856_out;
SharedReg704_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg704_out;
   MUX_Product325_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg680_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg842_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg110_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg706_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg856_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg704_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg838_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg816_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg575_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg682_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg799_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg491_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg801_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg802_out_to_MUX_Product325_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product325_0_impl_1_out);

   Delay1No273_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product325_0_impl_1_out,
                 Y => Delay1No273_out);

Delay1No274_out_to_Product325_4_impl_parent_implementedSystem_port_0_cast <= Delay1No274_out;
Delay1No275_out_to_Product325_4_impl_parent_implementedSystem_port_1_cast <= Delay1No275_out;
   Product325_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product325_4_impl_out,
                 X => Delay1No274_out_to_Product325_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No275_out_to_Product325_4_impl_parent_implementedSystem_port_1_cast);

SharedReg794_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg794_out;
SharedReg795_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg795_out;
SharedReg820_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg820_out;
SharedReg518_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg518_out;
SharedReg777_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg777_out;
SharedReg801_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg801_out;
SharedReg231_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg231_out;
SharedReg803_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg803_out;
SharedReg855_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg855_out;
SharedReg851_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg851_out;
SharedReg833_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg833_out;
SharedReg700_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg700_out;
SharedReg728_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg728_out;
SharedReg699_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg699_out;
   MUX_Product325_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg794_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg795_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg833_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg700_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg728_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg699_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg820_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg518_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg777_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg801_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg231_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg803_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg855_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg851_out_to_MUX_Product325_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product325_4_impl_0_out);

   Delay1No274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product325_4_impl_0_out,
                 Y => Delay1No274_out);

SharedReg699_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg699_out;
SharedReg595_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg595_out;
SharedReg702_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg702_out;
SharedReg799_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg799_out;
SharedReg519_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg519_out;
SharedReg274_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg274_out;
SharedReg802_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg802_out;
SharedReg130_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg130_out;
SharedReg730_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg730_out;
SharedReg771_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg771_out;
SharedReg768_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg768_out;
SharedReg841_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg841_out;
SharedReg842_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg842_out;
SharedReg838_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg838_out;
   MUX_Product325_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg699_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg595_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg768_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg841_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg842_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg838_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg702_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg799_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg519_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg274_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg802_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg130_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg730_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg771_out_to_MUX_Product325_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product325_4_impl_1_out);

   Delay1No275_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product325_4_impl_1_out,
                 Y => Delay1No275_out);

Delay1No276_out_to_Subtract26_0_impl_parent_implementedSystem_port_0_cast <= Delay1No276_out;
Delay1No277_out_to_Subtract26_0_impl_parent_implementedSystem_port_1_cast <= Delay1No277_out;
   Subtract26_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract26_0_impl_out,
                 X => Delay1No276_out_to_Subtract26_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No277_out_to_Subtract26_0_impl_parent_implementedSystem_port_1_cast);

SharedReg201_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg201_out;
SharedReg4_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg4_out;
SharedReg10_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg10_out;
SharedReg410_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg410_out;
SharedReg548_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg548_out;
SharedReg327_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg327_out;
SharedReg470_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg470_out;
SharedReg202_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg202_out;
SharedReg326_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg326_out;
SharedReg330_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg330_out;
SharedReg160_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg160_out;
SharedReg495_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg495_out;
SharedReg107_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg107_out;
SharedReg490_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg490_out;
   MUX_Subtract26_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg201_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg4_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg160_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg495_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg107_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg490_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg10_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg410_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg548_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg327_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg470_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg202_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg326_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg330_out_to_MUX_Subtract26_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract26_0_impl_0_out);

   Delay1No276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_0_impl_0_out,
                 Y => Delay1No276_out);

SharedReg133_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg133_out;
SharedReg20_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg20_out;
SharedReg26_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg26_out;
SharedReg470_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg470_out;
SharedReg490_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg490_out;
SharedReg546_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg546_out;
SharedReg632_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg632_out;
SharedReg136_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg136_out;
SharedReg490_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg490_out;
SharedReg546_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg546_out;
SharedReg132_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg132_out;
SharedReg326_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg326_out;
SharedReg63_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg63_out;
SharedReg549_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg549_out;
   MUX_Subtract26_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg133_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg20_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg132_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg326_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg63_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg549_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg26_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg470_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg490_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg546_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg632_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg136_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg490_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg546_out_to_MUX_Subtract26_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract26_0_impl_1_out);

   Delay1No277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_0_impl_1_out,
                 Y => Delay1No277_out);

Delay1No278_out_to_Subtract26_1_impl_parent_implementedSystem_port_0_cast <= Delay1No278_out;
Delay1No279_out_to_Subtract26_1_impl_parent_implementedSystem_port_1_cast <= Delay1No279_out;
   Subtract26_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract26_1_impl_out,
                 X => Delay1No278_out_to_Subtract26_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No279_out_to_Subtract26_1_impl_parent_implementedSystem_port_1_cast);

SharedReg502_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg502_out;
SharedReg112_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg112_out;
SharedReg497_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg497_out;
SharedReg209_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg209_out;
SharedReg4_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg4_out;
SharedReg10_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg10_out;
SharedReg414_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg414_out;
SharedReg553_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg553_out;
SharedReg334_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg334_out;
SharedReg454_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg454_out;
SharedReg210_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg210_out;
SharedReg333_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg333_out;
SharedReg337_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg337_out;
SharedReg168_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg168_out;
   MUX_Subtract26_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg502_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg112_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg210_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg333_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg337_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg168_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg497_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg209_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg4_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg10_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg414_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg553_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg334_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg454_out_to_MUX_Subtract26_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract26_1_impl_0_out);

   Delay1No278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_1_impl_0_out,
                 Y => Delay1No278_out);

SharedReg333_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg333_out;
SharedReg69_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg69_out;
SharedReg554_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg554_out;
SharedReg138_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg138_out;
SharedReg20_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg20_out;
SharedReg26_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg26_out;
SharedReg475_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg475_out;
SharedReg497_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg497_out;
SharedReg551_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg551_out;
SharedReg621_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg621_out;
SharedReg141_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg141_out;
SharedReg497_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg497_out;
SharedReg551_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg551_out;
SharedReg137_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg137_out;
   MUX_Subtract26_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg333_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg69_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg141_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg497_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg551_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg137_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg554_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg138_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg20_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg26_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg475_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg497_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg551_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg621_out_to_MUX_Subtract26_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract26_1_impl_1_out);

   Delay1No279_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_1_impl_1_out,
                 Y => Delay1No279_out);

Delay1No280_out_to_Subtract26_2_impl_parent_implementedSystem_port_0_cast <= Delay1No280_out;
Delay1No281_out_to_Subtract26_2_impl_parent_implementedSystem_port_1_cast <= Delay1No281_out;
   Subtract26_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract26_2_impl_out,
                 X => Delay1No280_out_to_Subtract26_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No281_out_to_Subtract26_2_impl_parent_implementedSystem_port_1_cast);

SharedReg340_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg340_out;
SharedReg344_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg344_out;
SharedReg176_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg176_out;
SharedReg509_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg509_out;
SharedReg117_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg117_out;
SharedReg504_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg504_out;
SharedReg217_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg217_out;
SharedReg4_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg4_out;
SharedReg10_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg10_out;
SharedReg418_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg418_out;
SharedReg558_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg558_out;
SharedReg341_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg341_out;
SharedReg479_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg479_out;
SharedReg218_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg218_out;
   MUX_Subtract26_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg340_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg344_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg558_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg341_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg479_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg218_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg176_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg509_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg117_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg504_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg217_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg4_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg10_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg418_out_to_MUX_Subtract26_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract26_2_impl_0_out);

   Delay1No280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_2_impl_0_out,
                 Y => Delay1No280_out);

SharedReg504_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg504_out;
SharedReg556_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg556_out;
SharedReg142_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg142_out;
SharedReg340_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg340_out;
SharedReg75_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg75_out;
SharedReg559_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg559_out;
SharedReg143_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg143_out;
SharedReg20_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg20_out;
SharedReg26_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg26_out;
SharedReg479_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg479_out;
SharedReg504_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg504_out;
SharedReg556_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg556_out;
SharedReg626_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg626_out;
SharedReg146_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg146_out;
   MUX_Subtract26_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg504_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg556_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg504_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg556_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg626_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg146_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg142_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg340_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg75_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg559_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg143_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg20_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg26_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg479_out_to_MUX_Subtract26_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract26_2_impl_1_out);

   Delay1No281_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_2_impl_1_out,
                 Y => Delay1No281_out);

Delay1No282_out_to_Subtract26_3_impl_parent_implementedSystem_port_0_cast <= Delay1No282_out;
Delay1No283_out_to_Subtract26_3_impl_parent_implementedSystem_port_1_cast <= Delay1No283_out;
   Subtract26_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract26_3_impl_out,
                 X => Delay1No282_out_to_Subtract26_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No283_out_to_Subtract26_3_impl_parent_implementedSystem_port_1_cast);

SharedReg348_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg348_out;
SharedReg461_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg461_out;
SharedReg226_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg226_out;
SharedReg347_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg347_out;
SharedReg351_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg351_out;
SharedReg184_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg184_out;
SharedReg516_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg516_out;
SharedReg122_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg122_out;
SharedReg511_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg511_out;
SharedReg225_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg225_out;
SharedReg4_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg4_out;
SharedReg10_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg10_out;
SharedReg422_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg422_out;
SharedReg563_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg563_out;
   MUX_Subtract26_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg348_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg461_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg4_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg10_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg422_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg563_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg226_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg347_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg351_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg184_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg516_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg122_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg511_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg225_out_to_MUX_Subtract26_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract26_3_impl_0_out);

   Delay1No282_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_3_impl_0_out,
                 Y => Delay1No282_out);

SharedReg561_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg561_out;
SharedReg605_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg605_out;
SharedReg151_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg151_out;
SharedReg511_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg511_out;
SharedReg561_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg561_out;
SharedReg147_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg147_out;
SharedReg347_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg347_out;
SharedReg81_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg81_out;
SharedReg564_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg564_out;
SharedReg148_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg148_out;
SharedReg20_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg20_out;
SharedReg26_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg26_out;
SharedReg482_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg482_out;
SharedReg511_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg511_out;
   MUX_Subtract26_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg561_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg605_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg20_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg26_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg482_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg511_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg151_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg511_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg561_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg147_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg347_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg81_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg564_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg148_out_to_MUX_Subtract26_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract26_3_impl_1_out);

   Delay1No283_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_3_impl_1_out,
                 Y => Delay1No283_out);

Delay1No284_out_to_Subtract26_4_impl_parent_implementedSystem_port_0_cast <= Delay1No284_out;
Delay1No285_out_to_Subtract26_4_impl_parent_implementedSystem_port_1_cast <= Delay1No285_out;
   Subtract26_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract26_4_impl_out,
                 X => Delay1No284_out_to_Subtract26_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No285_out_to_Subtract26_4_impl_parent_implementedSystem_port_1_cast);

SharedReg446_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg446_out;
SharedReg568_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg568_out;
SharedReg355_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg355_out;
SharedReg486_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg486_out;
SharedReg234_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg234_out;
SharedReg354_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg354_out;
SharedReg358_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg358_out;
SharedReg192_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg192_out;
SharedReg523_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg523_out;
SharedReg127_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg127_out;
SharedReg518_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg518_out;
SharedReg233_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg233_out;
SharedReg4_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg4_out;
SharedReg10_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg10_out;
   MUX_Subtract26_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg446_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg568_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg518_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg233_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg4_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg10_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg355_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg486_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg234_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg354_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg358_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg192_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg523_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg127_out_to_MUX_Subtract26_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract26_4_impl_0_out);

   Delay1No284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_4_impl_0_out,
                 Y => Delay1No284_out);

SharedReg542_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg542_out;
SharedReg518_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg518_out;
SharedReg566_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg566_out;
SharedReg635_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg635_out;
SharedReg156_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg156_out;
SharedReg518_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg518_out;
SharedReg566_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg566_out;
SharedReg152_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg152_out;
SharedReg354_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg354_out;
SharedReg87_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg87_out;
SharedReg569_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg569_out;
SharedReg153_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg153_out;
SharedReg20_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg20_out;
SharedReg26_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg26_out;
   MUX_Subtract26_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg542_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg518_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg569_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg153_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg20_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg26_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg566_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg635_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg156_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg518_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg566_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg152_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg354_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg87_out_to_MUX_Subtract26_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract26_4_impl_1_out);

   Delay1No285_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract26_4_impl_1_out,
                 Y => Delay1No285_out);

Delay1No286_out_to_Product55_1_impl_parent_implementedSystem_port_0_cast <= Delay1No286_out;
Delay1No287_out_to_Product55_1_impl_parent_implementedSystem_port_1_cast <= Delay1No287_out;
   Product55_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product55_1_impl_out,
                 X => Delay1No286_out_to_Product55_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No287_out_to_Product55_1_impl_parent_implementedSystem_port_1_cast);

SharedReg850_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg850_out;
SharedReg747_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg747_out;
SharedReg840_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg840_out;
SharedReg834_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg834_out;
SharedReg710_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg710_out;
SharedReg836_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg836_out;
SharedReg642_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg642_out;
SharedReg795_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg795_out;
SharedReg820_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg820_out;
SharedReg497_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg497_out;
SharedReg777_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg777_out;
SharedReg801_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg801_out;
SharedReg779_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg779_out;
SharedReg780_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg780_out;
   MUX_Product55_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg850_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg747_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg777_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg801_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg779_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg780_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg840_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg834_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg710_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg836_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg642_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg795_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg820_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg497_out_to_MUX_Product55_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product55_1_impl_0_out);

   Delay1No286_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_1_impl_0_out,
                 Y => Delay1No286_out);

SharedReg712_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg712_out;
SharedReg856_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg856_out;
SharedReg710_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg710_out;
SharedReg685_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg685_out;
SharedReg842_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg842_out;
SharedReg710_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg710_out;
SharedReg816_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg816_out;
SharedReg580_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg580_out;
SharedReg687_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg687_out;
SharedReg799_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg799_out;
SharedReg498_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg498_out;
SharedReg247_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg247_out;
SharedReg248_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg248_out;
SharedReg167_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg167_out;
   MUX_Product55_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg712_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg856_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg498_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg247_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg248_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg167_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg710_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg685_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg842_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg710_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg816_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg580_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg687_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg799_out_to_MUX_Product55_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product55_1_impl_1_out);

   Delay1No287_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_1_impl_1_out,
                 Y => Delay1No287_out);

Delay1No288_out_to_Product55_2_impl_parent_implementedSystem_port_0_cast <= Delay1No288_out;
Delay1No289_out_to_Product55_2_impl_parent_implementedSystem_port_1_cast <= Delay1No289_out;
   Product55_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product55_2_impl_out,
                 X => Delay1No288_out_to_Product55_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No289_out_to_Product55_2_impl_parent_implementedSystem_port_1_cast);

SharedReg801_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg801_out;
SharedReg779_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg779_out;
SharedReg780_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg780_out;
SharedReg850_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg850_out;
SharedReg755_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg755_out;
SharedReg752_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg752_out;
SharedReg834_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg834_out;
SharedReg716_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg716_out;
SharedReg836_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg836_out;
SharedReg647_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg647_out;
SharedReg795_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg795_out;
SharedReg647_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg647_out;
SharedReg862_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg862_out;
SharedReg863_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg863_out;
   MUX_Product55_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg801_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg779_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg795_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg647_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg862_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg863_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg780_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg850_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg755_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg752_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg834_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg716_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg836_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg647_out_to_MUX_Product55_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product55_2_impl_0_out);

   Delay1No288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_2_impl_0_out,
                 Y => Delay1No288_out);

SharedReg256_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg256_out;
SharedReg257_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg257_out;
SharedReg175_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg175_out;
SharedReg718_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg718_out;
SharedReg856_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg856_out;
SharedReg840_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg840_out;
SharedReg690_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg690_out;
SharedReg842_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg842_out;
SharedReg716_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg716_out;
SharedReg816_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg816_out;
SharedReg585_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg585_out;
SharedReg818_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg818_out;
SharedReg556_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg556_out;
SharedReg557_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg557_out;
   MUX_Product55_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg256_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg257_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg585_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg818_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg556_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg557_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg175_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg718_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg856_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg840_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg690_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg842_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg716_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg816_out_to_MUX_Product55_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product55_2_impl_1_out);

   Delay1No289_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_2_impl_1_out,
                 Y => Delay1No289_out);

Delay1No290_out_to_Product55_3_impl_parent_implementedSystem_port_0_cast <= Delay1No290_out;
Delay1No291_out_to_Product55_3_impl_parent_implementedSystem_port_1_cast <= Delay1No291_out;
   Product55_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product55_3_impl_out,
                 X => Delay1No290_out_to_Product55_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No291_out_to_Product55_3_impl_parent_implementedSystem_port_1_cast);

SharedReg652_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg652_out;
SharedReg862_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg862_out;
SharedReg863_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg863_out;
SharedReg801_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg801_out;
SharedReg779_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg779_out;
SharedReg803_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg803_out;
SharedReg850_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg850_out;
SharedReg763_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg763_out;
SharedReg760_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg760_out;
SharedReg834_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg834_out;
SharedReg722_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg722_out;
SharedReg843_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg843_out;
SharedReg794_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg794_out;
SharedReg795_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg795_out;
   MUX_Product55_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg652_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg862_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg722_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg843_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg794_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg795_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg863_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg801_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg779_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg803_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg850_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg763_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg760_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg834_out_to_MUX_Product55_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product55_3_impl_0_out);

   Delay1No290_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_3_impl_0_out,
                 Y => Delay1No290_out);

SharedReg818_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg818_out;
SharedReg561_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg561_out;
SharedReg562_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg562_out;
SharedReg265_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg265_out;
SharedReg266_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg266_out;
SharedReg183_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg183_out;
SharedReg724_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg724_out;
SharedReg856_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg856_out;
SharedReg840_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg840_out;
SharedReg695_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg695_out;
SharedReg842_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg842_out;
SharedReg722_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg722_out;
SharedReg694_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg694_out;
SharedReg762_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg762_out;
   MUX_Product55_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg818_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg561_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg842_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg722_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg694_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg762_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg562_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg265_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg266_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg183_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg724_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg856_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg840_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg695_out_to_MUX_Product55_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product55_3_impl_1_out);

   Delay1No291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product55_3_impl_1_out,
                 Y => Delay1No291_out);

Delay1No292_out_to_Product226_0_impl_parent_implementedSystem_port_0_cast <= Delay1No292_out;
Delay1No293_out_to_Product226_0_impl_parent_implementedSystem_port_1_cast <= Delay1No293_out;
   Product226_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product226_0_impl_out,
                 X => Delay1No292_out_to_Product226_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No293_out_to_Product226_0_impl_parent_implementedSystem_port_1_cast);

SharedReg680_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg680_out;
SharedReg835_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg835_out;
SharedReg836_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg836_out;
SharedReg794_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg794_out;
SharedReg795_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg795_out;
SharedReg637_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg637_out;
SharedReg862_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg862_out;
SharedReg863_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg863_out;
SharedReg801_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg801_out;
SharedReg779_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg779_out;
SharedReg780_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg780_out;
SharedReg855_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg855_out;
SharedReg781_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg781_out;
SharedReg736_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg736_out;
   MUX_Product226_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg680_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg835_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg780_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg855_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg781_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg736_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg836_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg794_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg795_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg637_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg862_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg863_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg801_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg779_out_to_MUX_Product226_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product226_0_impl_0_out);

   Delay1No292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_0_impl_0_out,
                 Y => Delay1No292_out);

SharedReg841_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg841_out;
SharedReg637_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg637_out;
SharedReg704_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg704_out;
SharedReg679_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg679_out;
SharedReg738_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg738_out;
SharedReg818_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg818_out;
SharedReg546_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg546_out;
SharedReg547_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg547_out;
SharedReg238_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg238_out;
SharedReg239_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg239_out;
SharedReg159_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg159_out;
SharedReg706_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg706_out;
SharedReg35_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg35_out;
SharedReg840_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg840_out;
   MUX_Product226_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg841_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg637_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg159_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg706_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg35_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg840_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg704_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg679_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg738_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg818_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg546_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg547_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg238_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg239_out_to_MUX_Product226_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product226_0_impl_1_out);

   Delay1No293_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_0_impl_1_out,
                 Y => Delay1No293_out);

Delay1No294_out_to_Product226_1_impl_parent_implementedSystem_port_0_cast <= Delay1No294_out;
Delay1No295_out_to_Product226_1_impl_parent_implementedSystem_port_1_cast <= Delay1No295_out;
   Product226_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product226_1_impl_out,
                 X => Delay1No294_out_to_Product226_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No295_out_to_Product226_1_impl_parent_implementedSystem_port_1_cast);

SharedReg855_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg855_out;
SharedReg781_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg781_out;
SharedReg744_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg744_out;
SharedReg685_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg685_out;
SharedReg835_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg835_out;
SharedReg843_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg843_out;
SharedReg794_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg794_out;
SharedReg795_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg795_out;
SharedReg642_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg642_out;
SharedReg862_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg862_out;
SharedReg863_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg863_out;
SharedReg248_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg248_out;
SharedReg779_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg779_out;
SharedReg803_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg803_out;
   MUX_Product226_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg855_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg781_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg863_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg248_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg779_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg803_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg744_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg685_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg835_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg843_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg794_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg795_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg642_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg862_out_to_MUX_Product226_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product226_1_impl_0_out);

   Delay1No294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_1_impl_0_out,
                 Y => Delay1No294_out);

SharedReg712_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg712_out;
SharedReg41_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg41_out;
SharedReg840_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg840_out;
SharedReg841_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg841_out;
SharedReg642_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg642_out;
SharedReg710_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg710_out;
SharedReg684_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg684_out;
SharedReg746_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg746_out;
SharedReg818_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg818_out;
SharedReg551_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg551_out;
SharedReg552_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg552_out;
SharedReg801_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg801_out;
SharedReg249_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg249_out;
SharedReg167_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg167_out;
   MUX_Product226_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg712_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg41_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg552_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg801_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg249_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg167_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg840_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg841_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg642_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg710_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg684_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg746_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg818_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg551_out_to_MUX_Product226_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Product226_1_impl_1_out);

   Delay1No295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product226_1_impl_1_out,
                 Y => Delay1No295_out);

Delay1No296_out_to_Product326_4_impl_parent_implementedSystem_port_0_cast <= Delay1No296_out;
Delay1No297_out_to_Product326_4_impl_parent_implementedSystem_port_1_cast <= Delay1No297_out;
   Product326_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product326_4_impl_out,
                 X => Delay1No296_out_to_Product326_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No297_out_to_Product326_4_impl_parent_implementedSystem_port_1_cast);

SharedReg275_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg275_out;
SharedReg771_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg771_out;
SharedReg657_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg657_out;
SharedReg699_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg699_out;
SharedReg836_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg836_out;
SharedReg835_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg835_out;
SharedReg840_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg840_out;
SharedReg795_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg795_out;
SharedReg780_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg780_out;
SharedReg804_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg804_out;
SharedReg779_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg779_out;
SharedReg862_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg862_out;
SharedReg863_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg863_out;
   MUX_Product326_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg275_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg771_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg779_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg862_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg863_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg657_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg699_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg836_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg835_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg840_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg795_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg780_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg804_out_to_MUX_Product326_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product326_4_impl_0_LUT_out,
                 oMux => MUX_Product326_4_impl_0_out);

   Delay1No296_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product326_4_impl_0_out,
                 Y => Delay1No296_out);

SharedReg191_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg191_out;
SharedReg61_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg61_out;
SharedReg275_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg275_out;
SharedReg566_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg566_out;
SharedReg567_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg567_out;
SharedReg728_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg728_out;
SharedReg770_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg770_out;
SharedReg657_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg657_out;
SharedReg728_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg728_out;
SharedReg856_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg856_out;
SharedReg818_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg818_out;
SharedReg816_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg816_out;
SharedReg801_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg801_out;
   MUX_Product326_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg191_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg61_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg818_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg816_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg801_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg275_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg566_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg567_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg728_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg770_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg657_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg728_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg856_out_to_MUX_Product326_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product326_4_impl_1_LUT_out,
                 oMux => MUX_Product326_4_impl_1_out);

   Delay1No297_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product326_4_impl_1_out,
                 Y => Delay1No297_out);

Delay1No298_out_to_Subtract29_0_impl_parent_implementedSystem_port_0_cast <= Delay1No298_out;
Delay1No299_out_to_Subtract29_0_impl_parent_implementedSystem_port_1_cast <= Delay1No299_out;
   Subtract29_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract29_0_impl_out,
                 X => Delay1No298_out_to_Subtract29_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No299_out_to_Subtract29_0_impl_parent_implementedSystem_port_1_cast);

SharedReg492_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg492_out;
SharedReg5_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg5_out;
SharedReg11_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg11_out;
SharedReg525_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg525_out;
SharedReg239_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg239_out;
SharedReg158_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg158_out;
SharedReg430_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg430_out;
SharedReg578_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg578_out;
SharedReg92_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg92_out;
SharedReg332_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg332_out;
SharedReg494_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg494_out;
SharedReg162_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg162_out;
SharedReg93_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg93_out;
SharedReg238_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg238_out;
   MUX_Subtract29_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg492_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg5_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg494_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg162_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg93_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg238_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg11_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg525_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg239_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg158_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg430_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg578_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg92_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg332_out_to_MUX_Subtract29_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract29_0_impl_0_out);

   Delay1No298_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract29_0_impl_0_out,
                 Y => Delay1No298_out);

SharedReg326_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg326_out;
SharedReg21_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg21_out;
SharedReg27_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg27_out;
SharedReg670_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg670_out;
SharedReg157_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg157_out;
SharedReg197_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg197_out;
SharedReg377_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg377_out;
SharedReg709_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg709_out;
SharedReg107_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg107_out;
SharedReg331_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg331_out;
SharedReg326_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg326_out;
SharedReg32_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg32_out;
SharedReg157_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg157_out;
SharedReg240_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg240_out;
   MUX_Subtract29_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg326_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg21_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg326_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg32_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg157_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg240_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg27_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg670_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg157_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg197_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg377_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg709_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg107_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg331_out_to_MUX_Subtract29_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract29_0_impl_1_out);

   Delay1No299_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract29_0_impl_1_out,
                 Y => Delay1No299_out);

Delay1No300_out_to_Subtract29_1_impl_parent_implementedSystem_port_0_cast <= Delay1No300_out;
Delay1No301_out_to_Subtract29_1_impl_parent_implementedSystem_port_1_cast <= Delay1No301_out;
   Subtract29_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract29_1_impl_out,
                 X => Delay1No300_out_to_Subtract29_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No301_out_to_Subtract29_1_impl_parent_implementedSystem_port_1_cast);

SharedReg170_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg170_out;
SharedReg96_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg96_out;
SharedReg247_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg247_out;
SharedReg499_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg499_out;
SharedReg5_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg5_out;
SharedReg11_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg11_out;
SharedReg529_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg529_out;
SharedReg248_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg248_out;
SharedReg166_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg166_out;
SharedReg414_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg414_out;
SharedReg583_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg583_out;
SharedReg95_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg95_out;
SharedReg339_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg339_out;
SharedReg501_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg501_out;
   MUX_Subtract29_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg170_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg96_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg583_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg95_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg339_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg501_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg247_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg499_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg5_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg11_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg529_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg248_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg166_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg414_out_to_MUX_Subtract29_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract29_1_impl_0_out);

   Delay1No300_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract29_1_impl_0_out,
                 Y => Delay1No300_out);

SharedReg38_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg38_out;
SharedReg165_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg165_out;
SharedReg249_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg249_out;
SharedReg333_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg333_out;
SharedReg21_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg21_out;
SharedReg27_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg27_out;
SharedReg673_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg673_out;
SharedReg165_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg165_out;
SharedReg205_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg205_out;
SharedReg380_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg380_out;
SharedReg715_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg715_out;
SharedReg112_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg112_out;
SharedReg338_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg338_out;
SharedReg333_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg333_out;
   MUX_Subtract29_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg38_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg165_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg715_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg112_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg338_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg333_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg249_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg333_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg21_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg27_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg673_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg165_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg205_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg380_out_to_MUX_Subtract29_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract29_1_impl_1_out);

   Delay1No301_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract29_1_impl_1_out,
                 Y => Delay1No301_out);

Delay1No302_out_to_Subtract29_2_impl_parent_implementedSystem_port_0_cast <= Delay1No302_out;
Delay1No303_out_to_Subtract29_2_impl_parent_implementedSystem_port_1_cast <= Delay1No303_out;
   Subtract29_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract29_2_impl_out,
                 X => Delay1No302_out_to_Subtract29_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No303_out_to_Subtract29_2_impl_parent_implementedSystem_port_1_cast);

SharedReg98_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg98_out;
SharedReg346_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg346_out;
SharedReg508_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg508_out;
SharedReg178_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg178_out;
SharedReg99_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg99_out;
SharedReg256_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg256_out;
SharedReg506_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg506_out;
SharedReg5_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg5_out;
SharedReg11_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg11_out;
SharedReg534_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg534_out;
SharedReg257_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg257_out;
SharedReg174_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg174_out;
SharedReg439_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg439_out;
SharedReg588_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg588_out;
   MUX_Subtract29_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg98_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg346_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg257_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg174_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg439_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg588_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg508_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg178_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg99_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg256_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg506_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg5_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg11_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg534_out_to_MUX_Subtract29_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract29_2_impl_0_out);

   Delay1No302_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract29_2_impl_0_out,
                 Y => Delay1No302_out);

SharedReg117_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg117_out;
SharedReg345_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg345_out;
SharedReg340_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg340_out;
SharedReg44_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg44_out;
SharedReg173_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg173_out;
SharedReg258_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg258_out;
SharedReg340_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg340_out;
SharedReg21_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg21_out;
SharedReg27_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg27_out;
SharedReg664_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg664_out;
SharedReg173_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg173_out;
SharedReg213_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg213_out;
SharedReg401_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg401_out;
SharedReg721_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg721_out;
   MUX_Subtract29_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg117_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg345_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg173_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg213_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg401_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg721_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg340_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg44_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg173_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg258_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg340_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg21_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg27_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg664_out_to_MUX_Subtract29_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract29_2_impl_1_out);

   Delay1No303_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract29_2_impl_1_out,
                 Y => Delay1No303_out);

Delay1No304_out_to_Subtract29_3_impl_parent_implementedSystem_port_0_cast <= Delay1No304_out;
Delay1No305_out_to_Subtract29_3_impl_parent_implementedSystem_port_1_cast <= Delay1No305_out;
   Subtract29_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract29_3_impl_out,
                 X => Delay1No304_out_to_Subtract29_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No305_out_to_Subtract29_3_impl_parent_implementedSystem_port_1_cast);

SharedReg182_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg182_out;
SharedReg422_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg422_out;
SharedReg593_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg593_out;
SharedReg101_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg101_out;
SharedReg353_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg353_out;
SharedReg515_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg515_out;
SharedReg186_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg186_out;
SharedReg102_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg102_out;
SharedReg265_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg265_out;
SharedReg513_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg513_out;
SharedReg5_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg5_out;
SharedReg11_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg11_out;
SharedReg538_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg538_out;
SharedReg266_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg266_out;
   MUX_Subtract29_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg182_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg422_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg5_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg11_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg538_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg266_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg593_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg101_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg353_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg515_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg186_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg102_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg265_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg513_out_to_MUX_Subtract29_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract29_3_impl_0_out);

   Delay1No304_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract29_3_impl_0_out,
                 Y => Delay1No304_out);

SharedReg221_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg221_out;
SharedReg404_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg404_out;
SharedReg727_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg727_out;
SharedReg122_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg122_out;
SharedReg352_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg352_out;
SharedReg347_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg347_out;
SharedReg50_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg50_out;
SharedReg181_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg181_out;
SharedReg267_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg267_out;
SharedReg347_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg347_out;
SharedReg21_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg21_out;
SharedReg27_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg27_out;
SharedReg667_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg667_out;
SharedReg181_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg181_out;
   MUX_Subtract29_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg221_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg404_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg21_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg27_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg667_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg181_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg727_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg122_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg352_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg347_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg50_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg181_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg267_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg347_out_to_MUX_Subtract29_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract29_3_impl_1_out);

   Delay1No305_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract29_3_impl_1_out,
                 Y => Delay1No305_out);

Delay1No306_out_to_Subtract29_4_impl_parent_implementedSystem_port_0_cast <= Delay1No306_out;
Delay1No307_out_to_Subtract29_4_impl_parent_implementedSystem_port_1_cast <= Delay1No307_out;
   Subtract29_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract29_4_impl_out,
                 X => Delay1No306_out_to_Subtract29_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No307_out_to_Subtract29_4_impl_parent_implementedSystem_port_1_cast);

SharedReg611_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg611_out;
SharedReg275_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg275_out;
SharedReg190_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg190_out;
SharedReg446_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg446_out;
SharedReg598_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg598_out;
SharedReg104_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg104_out;
SharedReg360_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg360_out;
SharedReg522_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg522_out;
SharedReg194_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg194_out;
SharedReg105_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg105_out;
SharedReg274_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg274_out;
SharedReg520_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg520_out;
SharedReg5_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg5_out;
SharedReg11_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg11_out;
   MUX_Subtract29_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg611_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg275_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg274_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg520_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg5_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg11_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg190_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg446_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg598_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg104_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg360_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg522_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg194_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg105_out_to_MUX_Subtract29_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract29_4_impl_0_out);

   Delay1No306_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract29_4_impl_0_out,
                 Y => Delay1No306_out);

SharedReg734_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg734_out;
SharedReg189_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg189_out;
SharedReg229_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg229_out;
SharedReg391_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg391_out;
SharedReg733_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg733_out;
SharedReg127_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg127_out;
SharedReg359_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg359_out;
SharedReg354_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg354_out;
SharedReg56_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg56_out;
SharedReg189_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg189_out;
SharedReg276_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg276_out;
SharedReg354_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg354_out;
SharedReg21_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg21_out;
SharedReg27_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg27_out;
   MUX_Subtract29_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg734_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg189_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg276_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg354_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg21_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg27_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg229_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg391_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg733_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg127_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg359_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg354_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg56_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg189_out_to_MUX_Subtract29_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract29_4_impl_1_out);

   Delay1No307_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract29_4_impl_1_out,
                 Y => Delay1No307_out);

Delay1No308_out_to_Subtract33_0_impl_parent_implementedSystem_port_0_cast <= Delay1No308_out;
Delay1No309_out_to_Subtract33_0_impl_parent_implementedSystem_port_1_cast <= Delay1No309_out;
   Subtract33_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract33_0_impl_out,
                 X => Delay1No308_out_to_Subtract33_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No309_out_to_Subtract33_0_impl_parent_implementedSystem_port_1_cast);

SharedReg547_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg547_out;
SharedReg13_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg13_out;
SharedReg12_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg12_out;
SharedReg576_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg576_out;
SharedReg326_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg326_out;
SharedReg328_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg328_out;
SharedReg471_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg471_out;
SharedReg244_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg244_out;
SharedReg546_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg546_out;
SharedReg495_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg495_out;
SharedReg158_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg158_out;
SharedReg329_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg329_out;
SharedReg546_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg546_out;
SharedReg574_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg574_out;
   MUX_Subtract33_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg547_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg13_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg158_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg329_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg546_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg574_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg12_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg576_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg326_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg328_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg471_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg244_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg546_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg495_out_to_MUX_Subtract33_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract33_0_impl_0_out);

   Delay1No308_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract33_0_impl_0_out,
                 Y => Delay1No308_out);

SharedReg641_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg641_out;
SharedReg29_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg29_out;
SharedReg28_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg28_out;
SharedReg490_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg490_out;
SharedReg547_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg547_out;
SharedReg574_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg574_out;
SharedReg633_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg633_out;
SharedReg164_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg164_out;
SharedReg574_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg574_out;
SharedReg683_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg683_out;
SharedReg157_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg157_out;
SharedReg574_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg574_out;
SharedReg493_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg493_out;
SharedReg682_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg682_out;
   MUX_Subtract33_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg641_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg29_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg157_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg574_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg493_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg682_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg28_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg490_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg547_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg574_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg633_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg164_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg574_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg683_out_to_MUX_Subtract33_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract33_0_impl_1_out);

   Delay1No309_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract33_0_impl_1_out,
                 Y => Delay1No309_out);

Delay1No310_out_to_Subtract33_1_impl_parent_implementedSystem_port_0_cast <= Delay1No310_out;
Delay1No311_out_to_Subtract33_1_impl_parent_implementedSystem_port_1_cast <= Delay1No311_out;
   Subtract33_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract33_1_impl_out,
                 X => Delay1No310_out_to_Subtract33_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No311_out_to_Subtract33_1_impl_parent_implementedSystem_port_1_cast);

SharedReg336_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg336_out;
SharedReg551_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg551_out;
SharedReg579_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg579_out;
SharedReg552_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg552_out;
SharedReg13_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg13_out;
SharedReg12_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg12_out;
SharedReg581_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg581_out;
SharedReg333_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg333_out;
SharedReg335_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg335_out;
SharedReg476_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg476_out;
SharedReg253_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg253_out;
SharedReg551_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg551_out;
SharedReg502_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg502_out;
SharedReg166_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg166_out;
   MUX_Subtract33_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg336_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg551_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg253_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg551_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg502_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg166_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg579_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg552_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg13_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg12_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg581_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg333_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg335_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg476_out_to_MUX_Subtract33_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract33_1_impl_0_out);

   Delay1No310_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract33_1_impl_0_out,
                 Y => Delay1No310_out);

SharedReg579_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg579_out;
SharedReg500_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg500_out;
SharedReg687_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg687_out;
SharedReg646_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg646_out;
SharedReg29_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg29_out;
SharedReg28_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg28_out;
SharedReg497_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg497_out;
SharedReg552_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg552_out;
SharedReg579_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg579_out;
SharedReg663_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg663_out;
SharedReg172_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg172_out;
SharedReg579_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg579_out;
SharedReg688_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg688_out;
SharedReg165_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg165_out;
   MUX_Subtract33_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg579_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg500_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg172_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg579_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg688_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg165_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg687_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg646_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg29_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg28_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg497_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg552_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg579_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg663_out_to_MUX_Subtract33_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract33_1_impl_1_out);

   Delay1No311_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract33_1_impl_1_out,
                 Y => Delay1No311_out);

Delay1No312_out_to_Subtract33_2_impl_parent_implementedSystem_port_0_cast <= Delay1No312_out;
Delay1No313_out_to_Subtract33_2_impl_parent_implementedSystem_port_1_cast <= Delay1No313_out;
   Subtract33_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract33_2_impl_out,
                 X => Delay1No312_out_to_Subtract33_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No313_out_to_Subtract33_2_impl_parent_implementedSystem_port_1_cast);

SharedReg556_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg556_out;
SharedReg509_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg509_out;
SharedReg174_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg174_out;
SharedReg343_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg343_out;
SharedReg556_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg556_out;
SharedReg584_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg584_out;
SharedReg557_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg557_out;
SharedReg13_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg13_out;
SharedReg12_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg12_out;
SharedReg586_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg586_out;
SharedReg340_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg340_out;
SharedReg342_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg342_out;
SharedReg535_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg535_out;
SharedReg262_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg262_out;
   MUX_Subtract33_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg556_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg509_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg340_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg342_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg535_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg262_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg174_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg343_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg556_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg584_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg557_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg13_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg12_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg586_out_to_MUX_Subtract33_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract33_2_impl_0_out);

   Delay1No312_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract33_2_impl_0_out,
                 Y => Delay1No312_out);

SharedReg584_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg584_out;
SharedReg693_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg693_out;
SharedReg173_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg173_out;
SharedReg584_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg584_out;
SharedReg507_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg507_out;
SharedReg692_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg692_out;
SharedReg651_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg651_out;
SharedReg29_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg29_out;
SharedReg28_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg28_out;
SharedReg504_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg504_out;
SharedReg557_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg557_out;
SharedReg584_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg584_out;
SharedReg665_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg665_out;
SharedReg180_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg180_out;
   MUX_Subtract33_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg584_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg693_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg557_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg584_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg665_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg180_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg173_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg584_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg507_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg692_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg651_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg29_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg28_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg504_out_to_MUX_Subtract33_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract33_2_impl_1_out);

   Delay1No313_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract33_2_impl_1_out,
                 Y => Delay1No313_out);

Delay1No314_out_to_Subtract33_3_impl_parent_implementedSystem_port_0_cast <= Delay1No314_out;
Delay1No315_out_to_Subtract33_3_impl_parent_implementedSystem_port_1_cast <= Delay1No315_out;
   Subtract33_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract33_3_impl_out,
                 X => Delay1No314_out_to_Subtract33_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No315_out_to_Subtract33_3_impl_parent_implementedSystem_port_1_cast);

SharedReg349_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg349_out;
SharedReg539_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg539_out;
SharedReg271_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg271_out;
SharedReg561_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg561_out;
SharedReg516_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg516_out;
SharedReg182_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg182_out;
SharedReg350_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg350_out;
SharedReg561_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg561_out;
SharedReg589_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg589_out;
SharedReg562_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg562_out;
SharedReg13_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg13_out;
SharedReg12_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg12_out;
SharedReg591_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg591_out;
SharedReg347_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg347_out;
   MUX_Subtract33_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg349_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg539_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg13_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg12_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg591_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg347_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg271_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg561_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg516_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg182_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg350_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg561_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg589_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg562_out_to_MUX_Subtract33_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract33_3_impl_0_out);

   Delay1No314_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract33_3_impl_0_out,
                 Y => Delay1No314_out);

SharedReg589_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg589_out;
SharedReg668_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg668_out;
SharedReg188_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg188_out;
SharedReg589_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg589_out;
SharedReg698_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg698_out;
SharedReg181_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg181_out;
SharedReg589_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg589_out;
SharedReg514_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg514_out;
SharedReg697_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg697_out;
SharedReg656_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg656_out;
SharedReg29_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg29_out;
SharedReg28_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg28_out;
SharedReg511_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg511_out;
SharedReg562_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg562_out;
   MUX_Subtract33_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg589_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg668_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg29_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg28_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg511_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg562_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg188_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg589_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg698_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg181_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg589_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg514_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg697_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg656_out_to_MUX_Subtract33_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract33_3_impl_1_out);

   Delay1No315_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract33_3_impl_1_out,
                 Y => Delay1No315_out);

Delay1No316_out_to_Subtract33_4_impl_parent_implementedSystem_port_0_cast <= Delay1No316_out;
Delay1No317_out_to_Subtract33_4_impl_parent_implementedSystem_port_1_cast <= Delay1No317_out;
   Subtract33_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract33_4_impl_out,
                 X => Delay1No316_out_to_Subtract33_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No317_out_to_Subtract33_4_impl_parent_implementedSystem_port_1_cast);

SharedReg596_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg596_out;
SharedReg354_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg354_out;
SharedReg356_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg356_out;
SharedReg487_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg487_out;
SharedReg280_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg280_out;
SharedReg566_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg566_out;
SharedReg523_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg523_out;
SharedReg190_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg190_out;
SharedReg357_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg357_out;
SharedReg566_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg566_out;
SharedReg594_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg594_out;
SharedReg567_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg567_out;
SharedReg13_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg13_out;
SharedReg12_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg12_out;
   MUX_Subtract33_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg596_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg354_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg594_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg567_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg13_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg12_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg356_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg487_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg280_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg566_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg523_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg190_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg357_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg566_out_to_MUX_Subtract33_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract33_4_impl_0_out);

   Delay1No316_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract33_4_impl_0_out,
                 Y => Delay1No316_out);

SharedReg518_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg518_out;
SharedReg567_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg567_out;
SharedReg594_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg594_out;
SharedReg636_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg636_out;
SharedReg196_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg196_out;
SharedReg594_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg594_out;
SharedReg703_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg703_out;
SharedReg189_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg189_out;
SharedReg594_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg594_out;
SharedReg521_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg521_out;
SharedReg702_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg702_out;
SharedReg661_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg661_out;
SharedReg29_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg29_out;
SharedReg28_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg28_out;
   MUX_Subtract33_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg518_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg567_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg702_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg661_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg29_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg28_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg594_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg636_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg196_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg594_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg703_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg189_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg594_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg521_out_to_MUX_Subtract33_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract33_4_impl_1_out);

   Delay1No317_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract33_4_impl_1_out,
                 Y => Delay1No317_out);

Delay1No318_out_to_Product237_4_impl_parent_implementedSystem_port_0_cast <= Delay1No318_out;
Delay1No319_out_to_Product237_4_impl_parent_implementedSystem_port_1_cast <= Delay1No319_out;
   Product237_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product237_4_impl_out,
                 X => Delay1No318_out_to_Product237_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No319_out_to_Product237_4_impl_parent_implementedSystem_port_1_cast);

SharedReg595_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg595_out;
SharedReg657_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg657_out;
SharedReg768_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg768_out;
SharedReg843_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg843_out;
SharedReg817_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg817_out;
SharedReg803_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg803_out;
SharedReg781_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg781_out;
SharedReg779_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg779_out;
SharedReg862_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg862_out;
   MUX_Product237_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg595_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg657_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg768_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg843_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg817_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg803_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg781_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg779_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg862_out_to_MUX_Product237_4_impl_0_parent_implementedSystem_port_9_cast,
                 iSel => MUX_Product237_4_impl_0_LUT_out,
                 oMux => MUX_Product237_4_impl_0_out);

   Delay1No318_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product237_4_impl_0_out,
                 Y => Delay1No318_out);

SharedReg191_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg191_out;
SharedReg59_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg59_out;
SharedReg276_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg276_out;
SharedReg594_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg594_out;
SharedReg770_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg770_out;
SharedReg728_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg728_out;
SharedReg842_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg842_out;
SharedReg840_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg840_out;
SharedReg863_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg863_out;
   MUX_Product237_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg191_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg59_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg276_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg594_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg770_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg728_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg842_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg840_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg863_out_to_MUX_Product237_4_impl_1_parent_implementedSystem_port_9_cast,
                 iSel => MUX_Product237_4_impl_1_LUT_out,
                 oMux => MUX_Product237_4_impl_1_out);

   Delay1No319_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product237_4_impl_1_out,
                 Y => Delay1No319_out);

Delay1No320_out_to_Subtract38_0_impl_parent_implementedSystem_port_0_cast <= Delay1No320_out;
Delay1No321_out_to_Subtract38_0_impl_parent_implementedSystem_port_1_cast <= Delay1No321_out;
   Subtract38_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract38_0_impl_out,
                 X => Delay1No320_out_to_Subtract38_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No321_out_to_Subtract38_0_impl_parent_implementedSystem_port_1_cast);

SharedReg198_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg198_out;
SharedReg15_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg15_out;
SharedReg14_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg14_out;
SharedReg198_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg198_out;
SharedReg132_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg132_out;
SharedReg134_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg134_out;
SharedReg670_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg670_out;
SharedReg135_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg135_out;
SharedReg132_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg132_out;
SharedReg162_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg162_out;
SharedReg495_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg495_out;
SharedReg546_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg546_out;
SharedReg197_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg197_out;
SharedReg237_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg237_out;
   MUX_Subtract38_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg198_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg495_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg546_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg197_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg237_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg14_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg198_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg132_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg134_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg670_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg135_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg132_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg162_out_to_MUX_Subtract38_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract38_0_impl_0_out);

   Delay1No320_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract38_0_impl_0_out,
                 Y => Delay1No320_out);

SharedReg243_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg243_out;
SharedReg31_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg31_out;
SharedReg30_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg30_out;
SharedReg197_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg197_out;
SharedReg238_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg238_out;
SharedReg237_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg237_out;
SharedReg287_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg287_out;
SharedReg161_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg161_out;
SharedReg197_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg197_out;
SharedReg111_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg111_out;
SharedReg743_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg743_out;
SharedReg637_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg637_out;
SharedReg199_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg199_out;
SharedReg241_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg241_out;
   MUX_Subtract38_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg243_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg31_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg743_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg637_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg199_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg241_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg30_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg197_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg238_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg237_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg287_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg161_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg197_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg111_out_to_MUX_Subtract38_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract38_0_impl_1_out);

   Delay1No321_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract38_0_impl_1_out,
                 Y => Delay1No321_out);

Delay1No322_out_to_Subtract38_1_impl_parent_implementedSystem_port_0_cast <= Delay1No322_out;
Delay1No323_out_to_Subtract38_1_impl_parent_implementedSystem_port_1_cast <= Delay1No323_out;
   Subtract38_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract38_1_impl_out,
                 X => Delay1No322_out_to_Subtract38_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No323_out_to_Subtract38_1_impl_parent_implementedSystem_port_1_cast);

SharedReg551_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg551_out;
SharedReg205_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg205_out;
SharedReg246_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg246_out;
SharedReg206_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg206_out;
SharedReg15_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg15_out;
SharedReg14_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg14_out;
SharedReg206_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg206_out;
SharedReg137_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg137_out;
SharedReg139_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg139_out;
SharedReg662_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg662_out;
SharedReg140_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg140_out;
SharedReg137_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg137_out;
SharedReg170_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg170_out;
SharedReg502_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg502_out;
   MUX_Subtract38_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg551_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg205_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg140_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg137_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg170_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg502_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg246_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg206_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg15_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg14_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg206_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg137_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg139_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg662_out_to_MUX_Subtract38_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract38_1_impl_0_out);

   Delay1No322_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract38_1_impl_0_out,
                 Y => Delay1No322_out);

SharedReg642_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg642_out;
SharedReg207_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg207_out;
SharedReg250_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg250_out;
SharedReg252_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg252_out;
SharedReg31_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg31_out;
SharedReg30_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg30_out;
SharedReg205_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg205_out;
SharedReg247_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg247_out;
SharedReg246_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg246_out;
SharedReg290_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg290_out;
SharedReg169_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg169_out;
SharedReg205_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg205_out;
SharedReg116_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg116_out;
SharedReg751_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg751_out;
   MUX_Subtract38_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg642_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg207_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg169_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg205_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg116_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg751_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg250_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg252_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg31_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg30_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg205_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg247_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg246_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg290_out_to_MUX_Subtract38_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract38_1_impl_1_out);

   Delay1No323_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract38_1_impl_1_out,
                 Y => Delay1No323_out);

Delay1No324_out_to_Subtract38_2_impl_parent_implementedSystem_port_0_cast <= Delay1No324_out;
Delay1No325_out_to_Subtract38_2_impl_parent_implementedSystem_port_1_cast <= Delay1No325_out;
   Subtract38_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract38_2_impl_out,
                 X => Delay1No324_out_to_Subtract38_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No325_out_to_Subtract38_2_impl_parent_implementedSystem_port_1_cast);

SharedReg142_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg142_out;
SharedReg178_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg178_out;
SharedReg509_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg509_out;
SharedReg556_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg556_out;
SharedReg213_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg213_out;
SharedReg255_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg255_out;
SharedReg214_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg214_out;
SharedReg15_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg15_out;
SharedReg14_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg14_out;
SharedReg214_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg214_out;
SharedReg142_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg142_out;
SharedReg144_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg144_out;
SharedReg664_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg664_out;
SharedReg145_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg145_out;
   MUX_Subtract38_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg142_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg178_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg142_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg144_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg664_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg145_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg509_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg556_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg213_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg255_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg214_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg15_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg14_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg214_out_to_MUX_Subtract38_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract38_2_impl_0_out);

   Delay1No324_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract38_2_impl_0_out,
                 Y => Delay1No324_out);

SharedReg213_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg213_out;
SharedReg121_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg121_out;
SharedReg759_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg759_out;
SharedReg647_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg647_out;
SharedReg215_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg215_out;
SharedReg259_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg259_out;
SharedReg261_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg261_out;
SharedReg31_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg31_out;
SharedReg30_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg30_out;
SharedReg213_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg213_out;
SharedReg256_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg256_out;
SharedReg255_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg255_out;
SharedReg293_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg293_out;
SharedReg177_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg177_out;
   MUX_Subtract38_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg213_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg121_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg256_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg255_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg293_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg177_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg759_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg647_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg215_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg259_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg261_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg31_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg30_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg213_out_to_MUX_Subtract38_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract38_2_impl_1_out);

   Delay1No325_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract38_2_impl_1_out,
                 Y => Delay1No325_out);

Delay1No326_out_to_Subtract38_3_impl_parent_implementedSystem_port_0_cast <= Delay1No326_out;
Delay1No327_out_to_Subtract38_3_impl_parent_implementedSystem_port_1_cast <= Delay1No327_out;
   Subtract38_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract38_3_impl_out,
                 X => Delay1No326_out_to_Subtract38_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No327_out_to_Subtract38_3_impl_parent_implementedSystem_port_1_cast);

SharedReg149_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg149_out;
SharedReg629_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg629_out;
SharedReg150_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg150_out;
SharedReg147_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg147_out;
SharedReg186_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg186_out;
SharedReg516_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg516_out;
SharedReg561_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg561_out;
SharedReg221_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg221_out;
SharedReg264_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg264_out;
SharedReg222_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg222_out;
SharedReg15_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg15_out;
SharedReg14_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg14_out;
SharedReg222_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg222_out;
SharedReg147_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg147_out;
   MUX_Subtract38_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg149_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg629_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg15_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg14_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg222_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg147_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg150_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg147_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg186_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg516_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg561_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg221_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg264_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg222_out_to_MUX_Subtract38_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract38_3_impl_0_out);

   Delay1No326_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract38_3_impl_0_out,
                 Y => Delay1No326_out);

SharedReg264_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg264_out;
SharedReg301_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg301_out;
SharedReg185_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg185_out;
SharedReg221_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg221_out;
SharedReg126_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg126_out;
SharedReg767_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg767_out;
SharedReg652_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg652_out;
SharedReg223_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg223_out;
SharedReg268_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg268_out;
SharedReg270_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg270_out;
SharedReg31_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg31_out;
SharedReg30_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg30_out;
SharedReg221_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg221_out;
SharedReg265_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg265_out;
   MUX_Subtract38_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg264_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg301_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg31_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg30_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg221_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg265_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg185_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg221_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg126_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg767_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg652_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg223_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg268_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg270_out_to_MUX_Subtract38_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract38_3_impl_1_out);

   Delay1No327_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract38_3_impl_1_out,
                 Y => Delay1No327_out);

Delay1No328_out_to_Subtract38_4_impl_parent_implementedSystem_port_0_cast <= Delay1No328_out;
Delay1No329_out_to_Subtract38_4_impl_parent_implementedSystem_port_1_cast <= Delay1No329_out;
   Subtract38_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract38_4_impl_out,
                 X => Delay1No328_out_to_Subtract38_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No329_out_to_Subtract38_4_impl_parent_implementedSystem_port_1_cast);

SharedReg230_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg230_out;
SharedReg152_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg152_out;
SharedReg154_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg154_out;
SharedReg676_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg676_out;
SharedReg155_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg155_out;
SharedReg152_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg152_out;
SharedReg194_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg194_out;
SharedReg523_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg523_out;
SharedReg566_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg566_out;
SharedReg229_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg229_out;
SharedReg273_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg273_out;
SharedReg230_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg230_out;
SharedReg15_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg15_out;
SharedReg14_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_14_cast <= SharedReg14_out;
   MUX_Subtract38_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg230_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg152_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg273_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg230_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg15_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg14_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg154_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg676_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg155_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg152_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg194_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg523_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg566_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg229_out_to_MUX_Subtract38_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract38_4_impl_0_out);

   Delay1No328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract38_4_impl_0_out,
                 Y => Delay1No328_out);

SharedReg229_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg229_out;
SharedReg274_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg274_out;
SharedReg273_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg273_out;
SharedReg735_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg735_out;
SharedReg193_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg193_out;
SharedReg229_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg229_out;
SharedReg131_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg131_out;
SharedReg775_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg775_out;
SharedReg657_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg657_out;
SharedReg231_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg231_out;
SharedReg277_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg277_out;
SharedReg279_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg279_out;
SharedReg31_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg31_out;
SharedReg30_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_14_cast <= SharedReg30_out;
   MUX_Subtract38_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_14_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg229_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg274_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg277_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg279_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg31_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg30_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_14_cast,
                 iS_2 => SharedReg273_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg735_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg193_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg229_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg131_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg775_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg657_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg231_out_to_MUX_Subtract38_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount141_out,
                 oMux => MUX_Subtract38_4_impl_1_out);

   Delay1No329_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract38_4_impl_1_out,
                 Y => Delay1No329_out);
   Constant2_0_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant2_0_impl_out);
   Constant11_0_impl_instance: Constant_float_8_23_0_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant11_0_impl_out);
   Constant4_0_impl_instance: Constant_float_8_23_cosnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant4_0_impl_out);
   Constant13_0_impl_instance: Constant_float_8_23_sinnpi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant13_0_impl_out);
   Constant5_0_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant5_0_impl_out);
   Constant14_0_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant14_0_impl_out);
   Constant6_0_impl_instance: Constant_float_8_23_cosnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant6_0_impl_out);
   Constant15_0_impl_instance: Constant_float_8_23_sinnpi_div_2_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant15_0_impl_out);
   Constant7_0_impl_instance: Constant_float_8_23_cosn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant7_0_impl_out);
   Constant16_0_impl_instance: Constant_float_8_23_sinn5_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant16_0_impl_out);
   Constant8_0_impl_instance: Constant_float_8_23_cosn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant8_0_impl_out);
   Constant17_0_impl_instance: Constant_float_8_23_sinn3_mult_pi_div_4_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant17_0_impl_out);
   Constant9_0_impl_instance: Constant_float_8_23_cosn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant9_0_impl_out);
   Constant18_0_impl_instance: Constant_float_8_23_sinn7_mult_pi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant18_0_impl_out);
   Constant_0_impl_instance: Constant_float_8_23_cosnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_0_impl_out);
   Constant1_0_impl_instance: Constant_float_8_23_sinnpi_div_8_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_0_impl_out);

   Delay9No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg37_out,
                 Y => Delay9No_out);

   Delay9No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => Delay9No1_out);

   Delay9No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => Delay9No2_out);

   Delay9No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg55_out,
                 Y => Delay9No3_out);

   Delay9No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => Delay9No4_out);

   Delay10No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => Delay10No_out);

   Delay10No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg73_out,
                 Y => Delay10No1_out);

   Delay10No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => Delay10No2_out);

   Delay10No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg85_out,
                 Y => Delay10No3_out);

   Delay10No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => Delay10No4_out);

   Delay10No25_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg528_out,
                 Y => Delay10No25_out);

   Delay10No26_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg533_out,
                 Y => Delay10No26_out);

   Delay10No27_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg537_out,
                 Y => Delay10No27_out);

   Delay10No28_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg541_out,
                 Y => Delay10No28_out);

   Delay10No29_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg545_out,
                 Y => Delay10No29_out);

   Delay4No71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg299_out,
                 Y => Delay4No71_out);

   Delay4No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg296_out,
                 Y => Delay4No74_out);

   Delay5No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg285_out,
                 Y => Delay5No10_out);

   Delay5No11_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg288_out,
                 Y => Delay5No11_out);

   Delay5No12_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg291_out,
                 Y => Delay5No12_out);

   Delay5No13_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg573_out,
                 Y => Delay5No13_out);

   Delay5No14_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg302_out,
                 Y => Delay5No14_out);

   Delay4No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg363_out,
                 Y => Delay4No75_out);

   Delay4No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg366_out,
                 Y => Delay4No76_out);

   Delay5No42_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg628_out,
                 Y => Delay5No42_out);

   Delay5No43_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg631_out,
                 Y => Delay5No43_out);

   Delay3No206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg663_out,
                 Y => Delay3No206_out);

   Delay3No214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg636_out,
                 Y => Delay3No214_out);

   Delay15No10_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg306_out,
                 Y => Delay15No10_out);

   Delay15No11_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg320_out,
                 Y => Delay15No11_out);

   Delay15No12_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg311_out,
                 Y => Delay15No12_out);

   Delay15No13_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg316_out,
                 Y => Delay15No13_out);

   Delay15No14_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg325_out,
                 Y => Delay15No14_out);

   Delay15No15_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg378_out,
                 Y => Delay15No15_out);

   Delay15No16_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg381_out,
                 Y => Delay15No16_out);

   Delay15No17_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg385_out,
                 Y => Delay15No17_out);

   Delay15No18_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg389_out,
                 Y => Delay15No18_out);

   Delay15No19_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg392_out,
                 Y => Delay15No19_out);

   Delay28No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => Delay28No_out);

   Delay28No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => Delay28No1_out);

   Delay28No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg121_out,
                 Y => Delay28No2_out);

   Delay28No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg126_out,
                 Y => Delay28No3_out);

   Delay28No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => Delay28No4_out);

   Delay15No20_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg395_out,
                 Y => Delay15No20_out);

   Delay15No21_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg399_out,
                 Y => Delay15No21_out);

   Delay15No22_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg402_out,
                 Y => Delay15No22_out);

   Delay15No23_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg406_out,
                 Y => Delay15No23_out);

   Delay15No24_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg409_out,
                 Y => Delay15No24_out);

   Delay15No25_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg413_out,
                 Y => Delay15No25_out);

   Delay15No26_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg417_out,
                 Y => Delay15No26_out);

   Delay15No27_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg421_out,
                 Y => Delay15No27_out);

   Delay15No28_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg425_out,
                 Y => Delay15No28_out);

   Delay15No29_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg429_out,
                 Y => Delay15No29_out);

   Delay15No30_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg434_out,
                 Y => Delay15No30_out);

   Delay15No31_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg438_out,
                 Y => Delay15No31_out);

   Delay15No32_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg442_out,
                 Y => Delay15No32_out);

   Delay15No33_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg445_out,
                 Y => Delay15No33_out);

   Delay15No34_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg449_out,
                 Y => Delay15No34_out);

   Delay15No35_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg453_out,
                 Y => Delay15No35_out);

   Delay15No36_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg456_out,
                 Y => Delay15No36_out);

   Delay15No37_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg460_out,
                 Y => Delay15No37_out);

   Delay15No38_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg465_out,
                 Y => Delay15No38_out);

   Delay15No39_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg469_out,
                 Y => Delay15No39_out);

   Delay10No60_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg578_out,
                 Y => Delay10No60_out);

   Delay10No61_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg583_out,
                 Y => Delay10No61_out);

   Delay10No62_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg588_out,
                 Y => Delay10No62_out);

   Delay10No63_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg593_out,
                 Y => Delay10No63_out);

   Delay10No64_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg598_out,
                 Y => Delay10No64_out);

   Delay27No15_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg164_out,
                 Y => Delay27No15_out);

   Delay27No16_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg172_out,
                 Y => Delay27No16_out);

   Delay27No17_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg180_out,
                 Y => Delay27No17_out);

   Delay27No18_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => Delay27No18_out);

   Delay27No19_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg196_out,
                 Y => Delay27No19_out);

   Delay27No20_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg709_out,
                 Y => Delay27No20_out);

   Delay27No21_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg715_out,
                 Y => Delay27No21_out);

   Delay27No22_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg721_out,
                 Y => Delay27No22_out);

   Delay27No23_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg727_out,
                 Y => Delay27No23_out);

   Delay27No24_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg733_out,
                 Y => Delay27No24_out);

   Delay16No_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg620_out,
                 Y => Delay16No_out);

   Delay16No1_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg625_out,
                 Y => Delay16No1_out);

   Delay16No2_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg604_out,
                 Y => Delay16No2_out);

   Delay16No3_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg610_out,
                 Y => Delay16No3_out);

   Delay16No4_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg615_out,
                 Y => Delay16No4_out);

   Delay16No5_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg672_out,
                 Y => Delay16No5_out);

   Delay16No6_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg675_out,
                 Y => Delay16No6_out);

   Delay16No7_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg666_out,
                 Y => Delay16No7_out);

   Delay16No8_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg669_out,
                 Y => Delay16No8_out);

   Delay16No9_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg678_out,
                 Y => Delay16No9_out);

   Delay3No249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg735_out,
                 Y => Delay3No249_out);

   Delay11No30_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg474_out,
                 Y => Delay11No30_out);

   Delay11No31_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg478_out,
                 Y => Delay11No31_out);

   Delay11No32_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg481_out,
                 Y => Delay11No32_out);

   Delay11No33_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg485_out,
                 Y => Delay11No33_out);

   Delay11No34_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg489_out,
                 Y => Delay11No34_out);

   Delay3No252_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg293_out,
                 Y => Delay3No252_out);

   MUX_y0_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y0_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y0_re_0_0_LUT_out);

   MUX_y0_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y0_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y0_im_0_0_LUT_out);

   MUX_y1_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y1_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y1_re_0_0_LUT_out);

   MUX_y1_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y1_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y1_im_0_0_LUT_out);

   MUX_y2_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y2_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y2_re_0_0_LUT_out);

   MUX_y2_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y2_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y2_im_0_0_LUT_out);

   MUX_y3_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y3_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y3_re_0_0_LUT_out);

   MUX_y3_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y3_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y3_im_0_0_LUT_out);

   MUX_y4_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y4_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y4_re_0_0_LUT_out);

   MUX_y4_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y4_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y4_im_0_0_LUT_out);

   MUX_y5_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y5_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y5_re_0_0_LUT_out);

   MUX_y5_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y5_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y5_im_0_0_LUT_out);

   MUX_y6_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y6_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y6_re_0_0_LUT_out);

   MUX_y6_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y6_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y6_im_0_0_LUT_out);

   MUX_y7_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y7_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y7_re_0_0_LUT_out);

   MUX_y7_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y7_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y7_im_0_0_LUT_out);

   MUX_y8_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y8_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y8_re_0_0_LUT_out);

   MUX_y8_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y8_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y8_im_0_0_LUT_out);

   MUX_y9_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y9_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y9_re_0_0_LUT_out);

   MUX_y9_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y9_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y9_im_0_0_LUT_out);

   MUX_y10_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y10_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y10_re_0_0_LUT_out);

   MUX_y10_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y10_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y10_im_0_0_LUT_out);

   MUX_y11_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y11_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y11_re_0_0_LUT_out);

   MUX_y11_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y11_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y11_im_0_0_LUT_out);

   MUX_y12_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y12_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y12_re_0_0_LUT_out);

   MUX_y12_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y12_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y12_im_0_0_LUT_out);

   MUX_y13_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y13_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y13_re_0_0_LUT_out);

   MUX_y13_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y13_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y13_im_0_0_LUT_out);

   MUX_y14_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y14_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y14_re_0_0_LUT_out);

   MUX_y14_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y14_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y14_im_0_0_LUT_out);

   MUX_y15_re_0_0_LUT_instance: GenericLut_LUTData_MUX_y15_re_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y15_re_0_0_LUT_out);

   MUX_y15_im_0_0_LUT_instance: GenericLut_LUTData_MUX_y15_im_0_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_y15_im_0_0_LUT_out);

   MUX_Product326_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product326_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Product326_4_impl_0_LUT_out);

   MUX_Product326_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product326_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Product326_4_impl_1_LUT_out);

   MUX_Product237_4_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product237_4_impl_0_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Product237_4_impl_0_LUT_out);

   MUX_Product237_4_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product237_4_impl_1_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount141_out,
                 Output => MUX_Product237_4_impl_1_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_re_0_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x0_im_0_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_re_0_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x1_im_0_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_re_0_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x2_im_0_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_re_0_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x3_im_0_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_re_0_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x4_im_0_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_re_0_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x5_im_0_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_re_0_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x6_im_0_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_re_0_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x7_im_0_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_re_0_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x8_im_0_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_re_0_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x9_im_0_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_re_0_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x10_im_0_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_re_0_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x11_im_0_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_re_0_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x12_im_0_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_re_0_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x13_im_0_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_re_0_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x14_im_0_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_re_0_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => x15_im_0_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_0_impl_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg33_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg34_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg35_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg36_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_1_impl_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg38_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg39_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg40_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_2_impl_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg47_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_3_impl_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add2_4_impl_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_0_impl_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg63_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_1_impl_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg69_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg71_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_2_impl_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg76_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_3_impl_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg80_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg81_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg82_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add11_4_impl_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg86_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg87_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg88_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg89_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg90_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_0_impl_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg92_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg93_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_1_impl_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg95_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_2_impl_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg98_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg99_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_3_impl_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg101_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg102_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add3_4_impl_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg104_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg105_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_0_impl_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg108_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg110_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_1_impl_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg112_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg113_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg115_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_2_impl_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg117_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg118_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_3_impl_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg123_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg125_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add12_4_impl_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg129_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add9_0_impl_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg132_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg134_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add9_1_impl_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg139_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg140_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add9_2_impl_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg143_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg144_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg145_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add9_3_impl_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add9_4_impl_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg152_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg153_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add18_0_impl_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg157_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg158_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg160_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg161_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg162_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg163_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add18_1_impl_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg166_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg167_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg168_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg169_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg170_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg171_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add18_2_impl_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg173_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg174_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg176_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg178_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg179_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add18_3_impl_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg181_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg182_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg183_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg184_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg185_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg186_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg187_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add18_4_impl_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg190_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg191_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg192_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg193_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg194_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg195_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add128_0_impl_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg197_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg198_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg200_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg201_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg202_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg203_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add128_1_impl_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg205_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg206_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg207_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg208_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg209_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg210_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg211_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add128_2_impl_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg213_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg214_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg215_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg216_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg217_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg218_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg219_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add128_3_impl_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg221_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg222_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg223_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg224_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg225_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg226_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg227_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add128_4_impl_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg229_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg230_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg231_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg232_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg233_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg234_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg235_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add40_0_impl_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg237_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg238_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg239_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg240_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg241_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg242_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg243_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg244_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add40_1_impl_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg246_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg247_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg248_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg250_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg251_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg252_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg253_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add40_2_impl_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg255_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg256_out,
                 Y => SharedReg257_out);

   SharedReg258_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg257_out,
                 Y => SharedReg258_out);

   SharedReg259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg258_out,
                 Y => SharedReg259_out);

   SharedReg260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg259_out,
                 Y => SharedReg260_out);

   SharedReg261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg260_out,
                 Y => SharedReg261_out);

   SharedReg262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg261_out,
                 Y => SharedReg262_out);

   SharedReg263_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg262_out,
                 Y => SharedReg263_out);

   SharedReg264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add40_3_impl_out,
                 Y => SharedReg264_out);

   SharedReg265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg264_out,
                 Y => SharedReg265_out);

   SharedReg266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg265_out,
                 Y => SharedReg266_out);

   SharedReg267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg266_out,
                 Y => SharedReg267_out);

   SharedReg268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg267_out,
                 Y => SharedReg268_out);

   SharedReg269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg268_out,
                 Y => SharedReg269_out);

   SharedReg270_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg269_out,
                 Y => SharedReg270_out);

   SharedReg271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg270_out,
                 Y => SharedReg271_out);

   SharedReg272_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg271_out,
                 Y => SharedReg272_out);

   SharedReg273_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add40_4_impl_out,
                 Y => SharedReg273_out);

   SharedReg274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg273_out,
                 Y => SharedReg274_out);

   SharedReg275_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg274_out,
                 Y => SharedReg275_out);

   SharedReg276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg275_out,
                 Y => SharedReg276_out);

   SharedReg277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg276_out,
                 Y => SharedReg277_out);

   SharedReg278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg277_out,
                 Y => SharedReg278_out);

   SharedReg279_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg278_out,
                 Y => SharedReg279_out);

   SharedReg280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg279_out,
                 Y => SharedReg280_out);

   SharedReg281_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg280_out,
                 Y => SharedReg281_out);

   SharedReg282_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_0_impl_out,
                 Y => SharedReg282_out);

   SharedReg283_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg282_out,
                 Y => SharedReg283_out);

   SharedReg284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg283_out,
                 Y => SharedReg284_out);

   SharedReg285_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg284_out,
                 Y => SharedReg285_out);

   SharedReg286_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_1_impl_out,
                 Y => SharedReg286_out);

   SharedReg287_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg286_out,
                 Y => SharedReg287_out);

   SharedReg288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg287_out,
                 Y => SharedReg288_out);

   SharedReg289_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_2_impl_out,
                 Y => SharedReg289_out);

   SharedReg290_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg289_out,
                 Y => SharedReg290_out);

   SharedReg291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg290_out,
                 Y => SharedReg291_out);

   SharedReg292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_3_impl_out,
                 Y => SharedReg292_out);

   SharedReg293_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg292_out,
                 Y => SharedReg293_out);

   SharedReg294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product4_4_impl_out,
                 Y => SharedReg294_out);

   SharedReg295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg294_out,
                 Y => SharedReg295_out);

   SharedReg296_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg295_out,
                 Y => SharedReg296_out);

   SharedReg297_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_1_impl_out,
                 Y => SharedReg297_out);

   SharedReg298_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg297_out,
                 Y => SharedReg298_out);

   SharedReg299_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg298_out,
                 Y => SharedReg299_out);

   SharedReg300_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product11_4_impl_out,
                 Y => SharedReg300_out);

   SharedReg301_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg300_out,
                 Y => SharedReg301_out);

   SharedReg302_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg301_out,
                 Y => SharedReg302_out);

   SharedReg303_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_0_impl_out,
                 Y => SharedReg303_out);

   SharedReg304_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg303_out,
                 Y => SharedReg304_out);

   SharedReg305_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg304_out,
                 Y => SharedReg305_out);

   SharedReg306_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg305_out,
                 Y => SharedReg306_out);

   SharedReg307_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_2_impl_out,
                 Y => SharedReg307_out);

   SharedReg308_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg307_out,
                 Y => SharedReg308_out);

   SharedReg309_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg308_out,
                 Y => SharedReg309_out);

   SharedReg310_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg309_out,
                 Y => SharedReg310_out);

   SharedReg311_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg310_out,
                 Y => SharedReg311_out);

   SharedReg312_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product21_3_impl_out,
                 Y => SharedReg312_out);

   SharedReg313_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg312_out,
                 Y => SharedReg313_out);

   SharedReg314_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg313_out,
                 Y => SharedReg314_out);

   SharedReg315_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg314_out,
                 Y => SharedReg315_out);

   SharedReg316_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg315_out,
                 Y => SharedReg316_out);

   SharedReg317_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_1_impl_out,
                 Y => SharedReg317_out);

   SharedReg318_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg317_out,
                 Y => SharedReg318_out);

   SharedReg319_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg318_out,
                 Y => SharedReg319_out);

   SharedReg320_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg319_out,
                 Y => SharedReg320_out);

   SharedReg321_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product31_4_impl_out,
                 Y => SharedReg321_out);

   SharedReg322_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg321_out,
                 Y => SharedReg322_out);

   SharedReg323_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg322_out,
                 Y => SharedReg323_out);

   SharedReg324_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg323_out,
                 Y => SharedReg324_out);

   SharedReg325_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg324_out,
                 Y => SharedReg325_out);

   SharedReg326_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_0_impl_out,
                 Y => SharedReg326_out);

   SharedReg327_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg326_out,
                 Y => SharedReg327_out);

   SharedReg328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg327_out,
                 Y => SharedReg328_out);

   SharedReg329_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg328_out,
                 Y => SharedReg329_out);

   SharedReg330_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg329_out,
                 Y => SharedReg330_out);

   SharedReg331_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg330_out,
                 Y => SharedReg331_out);

   SharedReg332_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg331_out,
                 Y => SharedReg332_out);

   SharedReg333_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_1_impl_out,
                 Y => SharedReg333_out);

   SharedReg334_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg333_out,
                 Y => SharedReg334_out);

   SharedReg335_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg334_out,
                 Y => SharedReg335_out);

   SharedReg336_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg335_out,
                 Y => SharedReg336_out);

   SharedReg337_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg336_out,
                 Y => SharedReg337_out);

   SharedReg338_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg337_out,
                 Y => SharedReg338_out);

   SharedReg339_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg338_out,
                 Y => SharedReg339_out);

   SharedReg340_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_2_impl_out,
                 Y => SharedReg340_out);

   SharedReg341_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg340_out,
                 Y => SharedReg341_out);

   SharedReg342_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg341_out,
                 Y => SharedReg342_out);

   SharedReg343_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg342_out,
                 Y => SharedReg343_out);

   SharedReg344_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg343_out,
                 Y => SharedReg344_out);

   SharedReg345_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg344_out,
                 Y => SharedReg345_out);

   SharedReg346_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg345_out,
                 Y => SharedReg346_out);

   SharedReg347_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_3_impl_out,
                 Y => SharedReg347_out);

   SharedReg348_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg347_out,
                 Y => SharedReg348_out);

   SharedReg349_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg348_out,
                 Y => SharedReg349_out);

   SharedReg350_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg349_out,
                 Y => SharedReg350_out);

   SharedReg351_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg350_out,
                 Y => SharedReg351_out);

   SharedReg352_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg351_out,
                 Y => SharedReg352_out);

   SharedReg353_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg352_out,
                 Y => SharedReg353_out);

   SharedReg354_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract2_4_impl_out,
                 Y => SharedReg354_out);

   SharedReg355_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg354_out,
                 Y => SharedReg355_out);

   SharedReg356_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg355_out,
                 Y => SharedReg356_out);

   SharedReg357_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg356_out,
                 Y => SharedReg357_out);

   SharedReg358_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg357_out,
                 Y => SharedReg358_out);

   SharedReg359_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg358_out,
                 Y => SharedReg359_out);

   SharedReg360_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg359_out,
                 Y => SharedReg360_out);

   SharedReg361_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product5_0_impl_out,
                 Y => SharedReg361_out);

   SharedReg362_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg361_out,
                 Y => SharedReg362_out);

   SharedReg363_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg362_out,
                 Y => SharedReg363_out);

   SharedReg364_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product5_1_impl_out,
                 Y => SharedReg364_out);

   SharedReg365_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg364_out,
                 Y => SharedReg365_out);

   SharedReg366_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg365_out,
                 Y => SharedReg366_out);

   SharedReg367_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product5_2_impl_out,
                 Y => SharedReg367_out);

   SharedReg368_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg367_out,
                 Y => SharedReg368_out);

   SharedReg369_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg368_out,
                 Y => SharedReg369_out);

   SharedReg370_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product5_3_impl_out,
                 Y => SharedReg370_out);

   SharedReg371_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg370_out,
                 Y => SharedReg371_out);

   SharedReg372_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg371_out,
                 Y => SharedReg372_out);

   SharedReg373_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product5_4_impl_out,
                 Y => SharedReg373_out);

   SharedReg374_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg373_out,
                 Y => SharedReg374_out);

   SharedReg375_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg374_out,
                 Y => SharedReg375_out);

   SharedReg376_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_0_impl_out,
                 Y => SharedReg376_out);

   SharedReg377_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg376_out,
                 Y => SharedReg377_out);

   SharedReg378_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg377_out,
                 Y => SharedReg378_out);

   SharedReg379_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_1_impl_out,
                 Y => SharedReg379_out);

   SharedReg380_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg379_out,
                 Y => SharedReg380_out);

   SharedReg381_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg380_out,
                 Y => SharedReg381_out);

   SharedReg382_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_2_impl_out,
                 Y => SharedReg382_out);

   SharedReg383_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg382_out,
                 Y => SharedReg383_out);

   SharedReg384_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg383_out,
                 Y => SharedReg384_out);

   SharedReg385_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg384_out,
                 Y => SharedReg385_out);

   SharedReg386_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_3_impl_out,
                 Y => SharedReg386_out);

   SharedReg387_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg386_out,
                 Y => SharedReg387_out);

   SharedReg388_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg387_out,
                 Y => SharedReg388_out);

   SharedReg389_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg388_out,
                 Y => SharedReg389_out);

   SharedReg390_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product12_4_impl_out,
                 Y => SharedReg390_out);

   SharedReg391_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg390_out,
                 Y => SharedReg391_out);

   SharedReg392_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg391_out,
                 Y => SharedReg392_out);

   SharedReg393_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_0_impl_out,
                 Y => SharedReg393_out);

   SharedReg394_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg393_out,
                 Y => SharedReg394_out);

   SharedReg395_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg394_out,
                 Y => SharedReg395_out);

   SharedReg396_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_1_impl_out,
                 Y => SharedReg396_out);

   SharedReg397_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg396_out,
                 Y => SharedReg397_out);

   SharedReg398_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg397_out,
                 Y => SharedReg398_out);

   SharedReg399_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg398_out,
                 Y => SharedReg399_out);

   SharedReg400_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_2_impl_out,
                 Y => SharedReg400_out);

   SharedReg401_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg400_out,
                 Y => SharedReg401_out);

   SharedReg402_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg401_out,
                 Y => SharedReg402_out);

   SharedReg403_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_3_impl_out,
                 Y => SharedReg403_out);

   SharedReg404_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg403_out,
                 Y => SharedReg404_out);

   SharedReg405_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg404_out,
                 Y => SharedReg405_out);

   SharedReg406_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg405_out,
                 Y => SharedReg406_out);

   SharedReg407_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product22_4_impl_out,
                 Y => SharedReg407_out);

   SharedReg408_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg407_out,
                 Y => SharedReg408_out);

   SharedReg409_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg408_out,
                 Y => SharedReg409_out);

   SharedReg410_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_0_impl_out,
                 Y => SharedReg410_out);

   SharedReg411_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg410_out,
                 Y => SharedReg411_out);

   SharedReg412_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg411_out,
                 Y => SharedReg412_out);

   SharedReg413_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg412_out,
                 Y => SharedReg413_out);

   SharedReg414_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_1_impl_out,
                 Y => SharedReg414_out);

   SharedReg415_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg414_out,
                 Y => SharedReg415_out);

   SharedReg416_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg415_out,
                 Y => SharedReg416_out);

   SharedReg417_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg416_out,
                 Y => SharedReg417_out);

   SharedReg418_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_2_impl_out,
                 Y => SharedReg418_out);

   SharedReg419_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg418_out,
                 Y => SharedReg419_out);

   SharedReg420_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg419_out,
                 Y => SharedReg420_out);

   SharedReg421_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg420_out,
                 Y => SharedReg421_out);

   SharedReg422_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_3_impl_out,
                 Y => SharedReg422_out);

   SharedReg423_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg422_out,
                 Y => SharedReg423_out);

   SharedReg424_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg423_out,
                 Y => SharedReg424_out);

   SharedReg425_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg424_out,
                 Y => SharedReg425_out);

   SharedReg426_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product32_4_impl_out,
                 Y => SharedReg426_out);

   SharedReg427_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg426_out,
                 Y => SharedReg427_out);

   SharedReg428_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg427_out,
                 Y => SharedReg428_out);

   SharedReg429_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg428_out,
                 Y => SharedReg429_out);

   SharedReg430_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_0_impl_out,
                 Y => SharedReg430_out);

   SharedReg431_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg430_out,
                 Y => SharedReg431_out);

   SharedReg432_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg431_out,
                 Y => SharedReg432_out);

   SharedReg433_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg432_out,
                 Y => SharedReg433_out);

   SharedReg434_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg433_out,
                 Y => SharedReg434_out);

   SharedReg435_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_1_impl_out,
                 Y => SharedReg435_out);

   SharedReg436_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg435_out,
                 Y => SharedReg436_out);

   SharedReg437_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg436_out,
                 Y => SharedReg437_out);

   SharedReg438_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg437_out,
                 Y => SharedReg438_out);

   SharedReg439_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_2_impl_out,
                 Y => SharedReg439_out);

   SharedReg440_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg439_out,
                 Y => SharedReg440_out);

   SharedReg441_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg440_out,
                 Y => SharedReg441_out);

   SharedReg442_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg441_out,
                 Y => SharedReg442_out);

   SharedReg443_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_3_impl_out,
                 Y => SharedReg443_out);

   SharedReg444_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg443_out,
                 Y => SharedReg444_out);

   SharedReg445_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg444_out,
                 Y => SharedReg445_out);

   SharedReg446_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product6_4_impl_out,
                 Y => SharedReg446_out);

   SharedReg447_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg446_out,
                 Y => SharedReg447_out);

   SharedReg448_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg447_out,
                 Y => SharedReg448_out);

   SharedReg449_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg448_out,
                 Y => SharedReg449_out);

   SharedReg450_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_0_impl_out,
                 Y => SharedReg450_out);

   SharedReg451_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg450_out,
                 Y => SharedReg451_out);

   SharedReg452_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg451_out,
                 Y => SharedReg452_out);

   SharedReg453_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg452_out,
                 Y => SharedReg453_out);

   SharedReg454_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_1_impl_out,
                 Y => SharedReg454_out);

   SharedReg455_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg454_out,
                 Y => SharedReg455_out);

   SharedReg456_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg455_out,
                 Y => SharedReg456_out);

   SharedReg457_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_2_impl_out,
                 Y => SharedReg457_out);

   SharedReg458_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg457_out,
                 Y => SharedReg458_out);

   SharedReg459_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg458_out,
                 Y => SharedReg459_out);

   SharedReg460_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg459_out,
                 Y => SharedReg460_out);

   SharedReg461_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_3_impl_out,
                 Y => SharedReg461_out);

   SharedReg462_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg461_out,
                 Y => SharedReg462_out);

   SharedReg463_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg462_out,
                 Y => SharedReg463_out);

   SharedReg464_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg463_out,
                 Y => SharedReg464_out);

   SharedReg465_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg464_out,
                 Y => SharedReg465_out);

   SharedReg466_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product23_4_impl_out,
                 Y => SharedReg466_out);

   SharedReg467_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg466_out,
                 Y => SharedReg467_out);

   SharedReg468_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg467_out,
                 Y => SharedReg468_out);

   SharedReg469_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg468_out,
                 Y => SharedReg469_out);

   SharedReg470_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_0_impl_out,
                 Y => SharedReg470_out);

   SharedReg471_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg470_out,
                 Y => SharedReg471_out);

   SharedReg472_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg471_out,
                 Y => SharedReg472_out);

   SharedReg473_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg472_out,
                 Y => SharedReg473_out);

   SharedReg474_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg473_out,
                 Y => SharedReg474_out);

   SharedReg475_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_1_impl_out,
                 Y => SharedReg475_out);

   SharedReg476_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg475_out,
                 Y => SharedReg476_out);

   SharedReg477_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg476_out,
                 Y => SharedReg477_out);

   SharedReg478_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg477_out,
                 Y => SharedReg478_out);

   SharedReg479_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_2_impl_out,
                 Y => SharedReg479_out);

   SharedReg480_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg479_out,
                 Y => SharedReg480_out);

   SharedReg481_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg480_out,
                 Y => SharedReg481_out);

   SharedReg482_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_3_impl_out,
                 Y => SharedReg482_out);

   SharedReg483_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg482_out,
                 Y => SharedReg483_out);

   SharedReg484_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg483_out,
                 Y => SharedReg484_out);

   SharedReg485_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg484_out,
                 Y => SharedReg485_out);

   SharedReg486_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product33_4_impl_out,
                 Y => SharedReg486_out);

   SharedReg487_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg486_out,
                 Y => SharedReg487_out);

   SharedReg488_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg487_out,
                 Y => SharedReg488_out);

   SharedReg489_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg488_out,
                 Y => SharedReg489_out);

   SharedReg490_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_0_impl_out,
                 Y => SharedReg490_out);

   SharedReg491_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg490_out,
                 Y => SharedReg491_out);

   SharedReg492_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg491_out,
                 Y => SharedReg492_out);

   SharedReg493_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg492_out,
                 Y => SharedReg493_out);

   SharedReg494_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg493_out,
                 Y => SharedReg494_out);

   SharedReg495_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg494_out,
                 Y => SharedReg495_out);

   SharedReg496_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg495_out,
                 Y => SharedReg496_out);

   SharedReg497_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_1_impl_out,
                 Y => SharedReg497_out);

   SharedReg498_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg497_out,
                 Y => SharedReg498_out);

   SharedReg499_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg498_out,
                 Y => SharedReg499_out);

   SharedReg500_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg499_out,
                 Y => SharedReg500_out);

   SharedReg501_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg500_out,
                 Y => SharedReg501_out);

   SharedReg502_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg501_out,
                 Y => SharedReg502_out);

   SharedReg503_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg502_out,
                 Y => SharedReg503_out);

   SharedReg504_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_2_impl_out,
                 Y => SharedReg504_out);

   SharedReg505_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg504_out,
                 Y => SharedReg505_out);

   SharedReg506_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg505_out,
                 Y => SharedReg506_out);

   SharedReg507_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg506_out,
                 Y => SharedReg507_out);

   SharedReg508_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg507_out,
                 Y => SharedReg508_out);

   SharedReg509_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg508_out,
                 Y => SharedReg509_out);

   SharedReg510_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg509_out,
                 Y => SharedReg510_out);

   SharedReg511_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_3_impl_out,
                 Y => SharedReg511_out);

   SharedReg512_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg511_out,
                 Y => SharedReg512_out);

   SharedReg513_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg512_out,
                 Y => SharedReg513_out);

   SharedReg514_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg513_out,
                 Y => SharedReg514_out);

   SharedReg515_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg514_out,
                 Y => SharedReg515_out);

   SharedReg516_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg515_out,
                 Y => SharedReg516_out);

   SharedReg517_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg516_out,
                 Y => SharedReg517_out);

   SharedReg518_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract4_4_impl_out,
                 Y => SharedReg518_out);

   SharedReg519_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg518_out,
                 Y => SharedReg519_out);

   SharedReg520_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg519_out,
                 Y => SharedReg520_out);

   SharedReg521_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg520_out,
                 Y => SharedReg521_out);

   SharedReg522_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg521_out,
                 Y => SharedReg522_out);

   SharedReg523_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg522_out,
                 Y => SharedReg523_out);

   SharedReg524_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg523_out,
                 Y => SharedReg524_out);

   SharedReg525_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product37_0_impl_out,
                 Y => SharedReg525_out);

   SharedReg526_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg525_out,
                 Y => SharedReg526_out);

   SharedReg527_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg526_out,
                 Y => SharedReg527_out);

   SharedReg528_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg527_out,
                 Y => SharedReg528_out);

   SharedReg529_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product37_1_impl_out,
                 Y => SharedReg529_out);

   SharedReg530_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg529_out,
                 Y => SharedReg530_out);

   SharedReg531_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg530_out,
                 Y => SharedReg531_out);

   SharedReg532_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg531_out,
                 Y => SharedReg532_out);

   SharedReg533_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg532_out,
                 Y => SharedReg533_out);

   SharedReg534_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product37_2_impl_out,
                 Y => SharedReg534_out);

   SharedReg535_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg534_out,
                 Y => SharedReg535_out);

   SharedReg536_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg535_out,
                 Y => SharedReg536_out);

   SharedReg537_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg536_out,
                 Y => SharedReg537_out);

   SharedReg538_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product37_3_impl_out,
                 Y => SharedReg538_out);

   SharedReg539_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg538_out,
                 Y => SharedReg539_out);

   SharedReg540_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg539_out,
                 Y => SharedReg540_out);

   SharedReg541_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg540_out,
                 Y => SharedReg541_out);

   SharedReg542_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product37_4_impl_out,
                 Y => SharedReg542_out);

   SharedReg543_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg542_out,
                 Y => SharedReg543_out);

   SharedReg544_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg543_out,
                 Y => SharedReg544_out);

   SharedReg545_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg544_out,
                 Y => SharedReg545_out);

   SharedReg546_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_0_impl_out,
                 Y => SharedReg546_out);

   SharedReg547_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg546_out,
                 Y => SharedReg547_out);

   SharedReg548_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg547_out,
                 Y => SharedReg548_out);

   SharedReg549_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg548_out,
                 Y => SharedReg549_out);

   SharedReg550_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg549_out,
                 Y => SharedReg550_out);

   SharedReg551_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_1_impl_out,
                 Y => SharedReg551_out);

   SharedReg552_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg551_out,
                 Y => SharedReg552_out);

   SharedReg553_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg552_out,
                 Y => SharedReg553_out);

   SharedReg554_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg553_out,
                 Y => SharedReg554_out);

   SharedReg555_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg554_out,
                 Y => SharedReg555_out);

   SharedReg556_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_2_impl_out,
                 Y => SharedReg556_out);

   SharedReg557_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg556_out,
                 Y => SharedReg557_out);

   SharedReg558_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg557_out,
                 Y => SharedReg558_out);

   SharedReg559_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg558_out,
                 Y => SharedReg559_out);

   SharedReg560_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg559_out,
                 Y => SharedReg560_out);

   SharedReg561_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_3_impl_out,
                 Y => SharedReg561_out);

   SharedReg562_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg561_out,
                 Y => SharedReg562_out);

   SharedReg563_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg562_out,
                 Y => SharedReg563_out);

   SharedReg564_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg563_out,
                 Y => SharedReg564_out);

   SharedReg565_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg564_out,
                 Y => SharedReg565_out);

   SharedReg566_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract9_4_impl_out,
                 Y => SharedReg566_out);

   SharedReg567_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg566_out,
                 Y => SharedReg567_out);

   SharedReg568_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg567_out,
                 Y => SharedReg568_out);

   SharedReg569_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg568_out,
                 Y => SharedReg569_out);

   SharedReg570_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg569_out,
                 Y => SharedReg570_out);

   SharedReg571_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product39_3_impl_out,
                 Y => SharedReg571_out);

   SharedReg572_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg571_out,
                 Y => SharedReg572_out);

   SharedReg573_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg572_out,
                 Y => SharedReg573_out);

   SharedReg574_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract20_0_impl_out,
                 Y => SharedReg574_out);

   SharedReg575_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg574_out,
                 Y => SharedReg575_out);

   SharedReg576_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg575_out,
                 Y => SharedReg576_out);

   SharedReg577_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg576_out,
                 Y => SharedReg577_out);

   SharedReg578_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg577_out,
                 Y => SharedReg578_out);

   SharedReg579_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract20_1_impl_out,
                 Y => SharedReg579_out);

   SharedReg580_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg579_out,
                 Y => SharedReg580_out);

   SharedReg581_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg580_out,
                 Y => SharedReg581_out);

   SharedReg582_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg581_out,
                 Y => SharedReg582_out);

   SharedReg583_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg582_out,
                 Y => SharedReg583_out);

   SharedReg584_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract20_2_impl_out,
                 Y => SharedReg584_out);

   SharedReg585_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg584_out,
                 Y => SharedReg585_out);

   SharedReg586_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg585_out,
                 Y => SharedReg586_out);

   SharedReg587_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg586_out,
                 Y => SharedReg587_out);

   SharedReg588_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg587_out,
                 Y => SharedReg588_out);

   SharedReg589_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract20_3_impl_out,
                 Y => SharedReg589_out);

   SharedReg590_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg589_out,
                 Y => SharedReg590_out);

   SharedReg591_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg590_out,
                 Y => SharedReg591_out);

   SharedReg592_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg591_out,
                 Y => SharedReg592_out);

   SharedReg593_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg592_out,
                 Y => SharedReg593_out);

   SharedReg594_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract20_4_impl_out,
                 Y => SharedReg594_out);

   SharedReg595_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg594_out,
                 Y => SharedReg595_out);

   SharedReg596_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg595_out,
                 Y => SharedReg596_out);

   SharedReg597_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg596_out,
                 Y => SharedReg597_out);

   SharedReg598_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg597_out,
                 Y => SharedReg598_out);

   SharedReg599_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product220_2_impl_out,
                 Y => SharedReg599_out);

   SharedReg600_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg599_out,
                 Y => SharedReg600_out);

   SharedReg601_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg600_out,
                 Y => SharedReg601_out);

   SharedReg602_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg601_out,
                 Y => SharedReg602_out);

   SharedReg603_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg602_out,
                 Y => SharedReg603_out);

   SharedReg604_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg603_out,
                 Y => SharedReg604_out);

   SharedReg605_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product220_3_impl_out,
                 Y => SharedReg605_out);

   SharedReg606_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg605_out,
                 Y => SharedReg606_out);

   SharedReg607_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg606_out,
                 Y => SharedReg607_out);

   SharedReg608_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg607_out,
                 Y => SharedReg608_out);

   SharedReg609_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg608_out,
                 Y => SharedReg609_out);

   SharedReg610_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg609_out,
                 Y => SharedReg610_out);

   SharedReg611_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product220_4_impl_out,
                 Y => SharedReg611_out);

   SharedReg612_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg611_out,
                 Y => SharedReg612_out);

   SharedReg613_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg612_out,
                 Y => SharedReg613_out);

   SharedReg614_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg613_out,
                 Y => SharedReg614_out);

   SharedReg615_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg614_out,
                 Y => SharedReg615_out);

   SharedReg616_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product323_0_impl_out,
                 Y => SharedReg616_out);

   SharedReg617_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg616_out,
                 Y => SharedReg617_out);

   SharedReg618_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg617_out,
                 Y => SharedReg618_out);

   SharedReg619_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg618_out,
                 Y => SharedReg619_out);

   SharedReg620_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg619_out,
                 Y => SharedReg620_out);

   SharedReg621_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product323_1_impl_out,
                 Y => SharedReg621_out);

   SharedReg622_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg621_out,
                 Y => SharedReg622_out);

   SharedReg623_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg622_out,
                 Y => SharedReg623_out);

   SharedReg624_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg623_out,
                 Y => SharedReg624_out);

   SharedReg625_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg624_out,
                 Y => SharedReg625_out);

   SharedReg626_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product323_2_impl_out,
                 Y => SharedReg626_out);

   SharedReg627_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg626_out,
                 Y => SharedReg627_out);

   SharedReg628_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg627_out,
                 Y => SharedReg628_out);

   SharedReg629_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product323_3_impl_out,
                 Y => SharedReg629_out);

   SharedReg630_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg629_out,
                 Y => SharedReg630_out);

   SharedReg631_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg630_out,
                 Y => SharedReg631_out);

   SharedReg632_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product325_0_impl_out,
                 Y => SharedReg632_out);

   SharedReg633_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg632_out,
                 Y => SharedReg633_out);

   SharedReg634_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg633_out,
                 Y => SharedReg634_out);

   SharedReg635_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product325_4_impl_out,
                 Y => SharedReg635_out);

   SharedReg636_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg635_out,
                 Y => SharedReg636_out);

   SharedReg637_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract26_0_impl_out,
                 Y => SharedReg637_out);

   SharedReg638_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg637_out,
                 Y => SharedReg638_out);

   SharedReg639_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg638_out,
                 Y => SharedReg639_out);

   SharedReg640_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg639_out,
                 Y => SharedReg640_out);

   SharedReg641_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg640_out,
                 Y => SharedReg641_out);

   SharedReg642_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract26_1_impl_out,
                 Y => SharedReg642_out);

   SharedReg643_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg642_out,
                 Y => SharedReg643_out);

   SharedReg644_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg643_out,
                 Y => SharedReg644_out);

   SharedReg645_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg644_out,
                 Y => SharedReg645_out);

   SharedReg646_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg645_out,
                 Y => SharedReg646_out);

   SharedReg647_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract26_2_impl_out,
                 Y => SharedReg647_out);

   SharedReg648_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg647_out,
                 Y => SharedReg648_out);

   SharedReg649_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg648_out,
                 Y => SharedReg649_out);

   SharedReg650_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg649_out,
                 Y => SharedReg650_out);

   SharedReg651_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg650_out,
                 Y => SharedReg651_out);

   SharedReg652_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract26_3_impl_out,
                 Y => SharedReg652_out);

   SharedReg653_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg652_out,
                 Y => SharedReg653_out);

   SharedReg654_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg653_out,
                 Y => SharedReg654_out);

   SharedReg655_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg654_out,
                 Y => SharedReg655_out);

   SharedReg656_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg655_out,
                 Y => SharedReg656_out);

   SharedReg657_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract26_4_impl_out,
                 Y => SharedReg657_out);

   SharedReg658_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg657_out,
                 Y => SharedReg658_out);

   SharedReg659_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg658_out,
                 Y => SharedReg659_out);

   SharedReg660_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg659_out,
                 Y => SharedReg660_out);

   SharedReg661_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg660_out,
                 Y => SharedReg661_out);

   SharedReg662_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product55_1_impl_out,
                 Y => SharedReg662_out);

   SharedReg663_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg662_out,
                 Y => SharedReg663_out);

   SharedReg664_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product55_2_impl_out,
                 Y => SharedReg664_out);

   SharedReg665_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg664_out,
                 Y => SharedReg665_out);

   SharedReg666_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg665_out,
                 Y => SharedReg666_out);

   SharedReg667_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product55_3_impl_out,
                 Y => SharedReg667_out);

   SharedReg668_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg667_out,
                 Y => SharedReg668_out);

   SharedReg669_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg668_out,
                 Y => SharedReg669_out);

   SharedReg670_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product226_0_impl_out,
                 Y => SharedReg670_out);

   SharedReg671_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg670_out,
                 Y => SharedReg671_out);

   SharedReg672_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg671_out,
                 Y => SharedReg672_out);

   SharedReg673_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product226_1_impl_out,
                 Y => SharedReg673_out);

   SharedReg674_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg673_out,
                 Y => SharedReg674_out);

   SharedReg675_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg674_out,
                 Y => SharedReg675_out);

   SharedReg676_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product326_4_impl_out,
                 Y => SharedReg676_out);

   SharedReg677_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg676_out,
                 Y => SharedReg677_out);

   SharedReg678_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg677_out,
                 Y => SharedReg678_out);

   SharedReg679_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract29_0_impl_out,
                 Y => SharedReg679_out);

   SharedReg680_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg679_out,
                 Y => SharedReg680_out);

   SharedReg681_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg680_out,
                 Y => SharedReg681_out);

   SharedReg682_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg681_out,
                 Y => SharedReg682_out);

   SharedReg683_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg682_out,
                 Y => SharedReg683_out);

   SharedReg684_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract29_1_impl_out,
                 Y => SharedReg684_out);

   SharedReg685_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg684_out,
                 Y => SharedReg685_out);

   SharedReg686_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg685_out,
                 Y => SharedReg686_out);

   SharedReg687_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg686_out,
                 Y => SharedReg687_out);

   SharedReg688_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg687_out,
                 Y => SharedReg688_out);

   SharedReg689_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract29_2_impl_out,
                 Y => SharedReg689_out);

   SharedReg690_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg689_out,
                 Y => SharedReg690_out);

   SharedReg691_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg690_out,
                 Y => SharedReg691_out);

   SharedReg692_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg691_out,
                 Y => SharedReg692_out);

   SharedReg693_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg692_out,
                 Y => SharedReg693_out);

   SharedReg694_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract29_3_impl_out,
                 Y => SharedReg694_out);

   SharedReg695_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg694_out,
                 Y => SharedReg695_out);

   SharedReg696_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg695_out,
                 Y => SharedReg696_out);

   SharedReg697_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg696_out,
                 Y => SharedReg697_out);

   SharedReg698_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg697_out,
                 Y => SharedReg698_out);

   SharedReg699_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract29_4_impl_out,
                 Y => SharedReg699_out);

   SharedReg700_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg699_out,
                 Y => SharedReg700_out);

   SharedReg701_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg700_out,
                 Y => SharedReg701_out);

   SharedReg702_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg701_out,
                 Y => SharedReg702_out);

   SharedReg703_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg702_out,
                 Y => SharedReg703_out);

   SharedReg704_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract33_0_impl_out,
                 Y => SharedReg704_out);

   SharedReg705_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg704_out,
                 Y => SharedReg705_out);

   SharedReg706_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg705_out,
                 Y => SharedReg706_out);

   SharedReg707_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg706_out,
                 Y => SharedReg707_out);

   SharedReg708_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg707_out,
                 Y => SharedReg708_out);

   SharedReg709_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg708_out,
                 Y => SharedReg709_out);

   SharedReg710_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract33_1_impl_out,
                 Y => SharedReg710_out);

   SharedReg711_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg710_out,
                 Y => SharedReg711_out);

   SharedReg712_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg711_out,
                 Y => SharedReg712_out);

   SharedReg713_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg712_out,
                 Y => SharedReg713_out);

   SharedReg714_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg713_out,
                 Y => SharedReg714_out);

   SharedReg715_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg714_out,
                 Y => SharedReg715_out);

   SharedReg716_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract33_2_impl_out,
                 Y => SharedReg716_out);

   SharedReg717_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg716_out,
                 Y => SharedReg717_out);

   SharedReg718_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg717_out,
                 Y => SharedReg718_out);

   SharedReg719_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg718_out,
                 Y => SharedReg719_out);

   SharedReg720_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg719_out,
                 Y => SharedReg720_out);

   SharedReg721_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg720_out,
                 Y => SharedReg721_out);

   SharedReg722_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract33_3_impl_out,
                 Y => SharedReg722_out);

   SharedReg723_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg722_out,
                 Y => SharedReg723_out);

   SharedReg724_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg723_out,
                 Y => SharedReg724_out);

   SharedReg725_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg724_out,
                 Y => SharedReg725_out);

   SharedReg726_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg725_out,
                 Y => SharedReg726_out);

   SharedReg727_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg726_out,
                 Y => SharedReg727_out);

   SharedReg728_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract33_4_impl_out,
                 Y => SharedReg728_out);

   SharedReg729_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg728_out,
                 Y => SharedReg729_out);

   SharedReg730_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg729_out,
                 Y => SharedReg730_out);

   SharedReg731_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg730_out,
                 Y => SharedReg731_out);

   SharedReg732_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg731_out,
                 Y => SharedReg732_out);

   SharedReg733_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg732_out,
                 Y => SharedReg733_out);

   SharedReg734_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product237_4_impl_out,
                 Y => SharedReg734_out);

   SharedReg735_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg734_out,
                 Y => SharedReg735_out);

   SharedReg736_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract38_0_impl_out,
                 Y => SharedReg736_out);

   SharedReg737_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg736_out,
                 Y => SharedReg737_out);

   SharedReg738_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg737_out,
                 Y => SharedReg738_out);

   SharedReg739_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg738_out,
                 Y => SharedReg739_out);

   SharedReg740_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg739_out,
                 Y => SharedReg740_out);

   SharedReg741_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg740_out,
                 Y => SharedReg741_out);

   SharedReg742_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg741_out,
                 Y => SharedReg742_out);

   SharedReg743_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg742_out,
                 Y => SharedReg743_out);

   SharedReg744_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract38_1_impl_out,
                 Y => SharedReg744_out);

   SharedReg745_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg744_out,
                 Y => SharedReg745_out);

   SharedReg746_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg745_out,
                 Y => SharedReg746_out);

   SharedReg747_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg746_out,
                 Y => SharedReg747_out);

   SharedReg748_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg747_out,
                 Y => SharedReg748_out);

   SharedReg749_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg748_out,
                 Y => SharedReg749_out);

   SharedReg750_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg749_out,
                 Y => SharedReg750_out);

   SharedReg751_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg750_out,
                 Y => SharedReg751_out);

   SharedReg752_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract38_2_impl_out,
                 Y => SharedReg752_out);

   SharedReg753_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg752_out,
                 Y => SharedReg753_out);

   SharedReg754_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg753_out,
                 Y => SharedReg754_out);

   SharedReg755_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg754_out,
                 Y => SharedReg755_out);

   SharedReg756_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg755_out,
                 Y => SharedReg756_out);

   SharedReg757_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg756_out,
                 Y => SharedReg757_out);

   SharedReg758_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg757_out,
                 Y => SharedReg758_out);

   SharedReg759_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg758_out,
                 Y => SharedReg759_out);

   SharedReg760_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract38_3_impl_out,
                 Y => SharedReg760_out);

   SharedReg761_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg760_out,
                 Y => SharedReg761_out);

   SharedReg762_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg761_out,
                 Y => SharedReg762_out);

   SharedReg763_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg762_out,
                 Y => SharedReg763_out);

   SharedReg764_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg763_out,
                 Y => SharedReg764_out);

   SharedReg765_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg764_out,
                 Y => SharedReg765_out);

   SharedReg766_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg765_out,
                 Y => SharedReg766_out);

   SharedReg767_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg766_out,
                 Y => SharedReg767_out);

   SharedReg768_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract38_4_impl_out,
                 Y => SharedReg768_out);

   SharedReg769_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg768_out,
                 Y => SharedReg769_out);

   SharedReg770_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg769_out,
                 Y => SharedReg770_out);

   SharedReg771_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg770_out,
                 Y => SharedReg771_out);

   SharedReg772_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg771_out,
                 Y => SharedReg772_out);

   SharedReg773_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg772_out,
                 Y => SharedReg773_out);

   SharedReg774_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg773_out,
                 Y => SharedReg774_out);

   SharedReg775_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg774_out,
                 Y => SharedReg775_out);

   SharedReg776_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant2_0_impl_out,
                 Y => SharedReg776_out);

   SharedReg777_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg776_out,
                 Y => SharedReg777_out);

   SharedReg778_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg777_out,
                 Y => SharedReg778_out);

   SharedReg779_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg778_out,
                 Y => SharedReg779_out);

   SharedReg780_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg779_out,
                 Y => SharedReg780_out);

   SharedReg781_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg780_out,
                 Y => SharedReg781_out);

   SharedReg782_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg781_out,
                 Y => SharedReg782_out);

   SharedReg783_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg782_out,
                 Y => SharedReg783_out);

   SharedReg784_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg783_out,
                 Y => SharedReg784_out);

   SharedReg785_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg784_out,
                 Y => SharedReg785_out);

   SharedReg786_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg785_out,
                 Y => SharedReg786_out);

   SharedReg787_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg786_out,
                 Y => SharedReg787_out);

   SharedReg788_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg787_out,
                 Y => SharedReg788_out);

   SharedReg789_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg788_out,
                 Y => SharedReg789_out);

   SharedReg790_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg789_out,
                 Y => SharedReg790_out);

   SharedReg791_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg790_out,
                 Y => SharedReg791_out);

   SharedReg792_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg791_out,
                 Y => SharedReg792_out);

   SharedReg793_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg792_out,
                 Y => SharedReg793_out);

   SharedReg794_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg793_out,
                 Y => SharedReg794_out);

   SharedReg795_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg794_out,
                 Y => SharedReg795_out);

   SharedReg796_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg795_out,
                 Y => SharedReg796_out);

   SharedReg797_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg796_out,
                 Y => SharedReg797_out);

   SharedReg798_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg797_out,
                 Y => SharedReg798_out);

   SharedReg799_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant11_0_impl_out,
                 Y => SharedReg799_out);

   SharedReg800_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg799_out,
                 Y => SharedReg800_out);

   SharedReg801_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg800_out,
                 Y => SharedReg801_out);

   SharedReg802_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg801_out,
                 Y => SharedReg802_out);

   SharedReg803_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg802_out,
                 Y => SharedReg803_out);

   SharedReg804_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg803_out,
                 Y => SharedReg804_out);

   SharedReg805_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg804_out,
                 Y => SharedReg805_out);

   SharedReg806_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg805_out,
                 Y => SharedReg806_out);

   SharedReg807_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg806_out,
                 Y => SharedReg807_out);

   SharedReg808_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg807_out,
                 Y => SharedReg808_out);

   SharedReg809_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg808_out,
                 Y => SharedReg809_out);

   SharedReg810_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg809_out,
                 Y => SharedReg810_out);

   SharedReg811_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg810_out,
                 Y => SharedReg811_out);

   SharedReg812_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg811_out,
                 Y => SharedReg812_out);

   SharedReg813_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg812_out,
                 Y => SharedReg813_out);

   SharedReg814_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg813_out,
                 Y => SharedReg814_out);

   SharedReg815_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg814_out,
                 Y => SharedReg815_out);

   SharedReg816_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg815_out,
                 Y => SharedReg816_out);

   SharedReg817_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg816_out,
                 Y => SharedReg817_out);

   SharedReg818_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg817_out,
                 Y => SharedReg818_out);

   SharedReg819_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg818_out,
                 Y => SharedReg819_out);

   SharedReg820_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg819_out,
                 Y => SharedReg820_out);

   SharedReg821_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant4_0_impl_out,
                 Y => SharedReg821_out);

   SharedReg822_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg821_out,
                 Y => SharedReg822_out);

   SharedReg823_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg822_out,
                 Y => SharedReg823_out);

   SharedReg824_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg823_out,
                 Y => SharedReg824_out);

   SharedReg825_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant13_0_impl_out,
                 Y => SharedReg825_out);

   SharedReg826_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg825_out,
                 Y => SharedReg826_out);

   SharedReg827_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg826_out,
                 Y => SharedReg827_out);

   SharedReg828_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant5_0_impl_out,
                 Y => SharedReg828_out);

   SharedReg829_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant14_0_impl_out,
                 Y => SharedReg829_out);

   SharedReg830_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant6_0_impl_out,
                 Y => SharedReg830_out);

   SharedReg831_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg830_out,
                 Y => SharedReg831_out);

   SharedReg832_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg831_out,
                 Y => SharedReg832_out);

   SharedReg833_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg832_out,
                 Y => SharedReg833_out);

   SharedReg834_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg833_out,
                 Y => SharedReg834_out);

   SharedReg835_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg834_out,
                 Y => SharedReg835_out);

   SharedReg836_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg835_out,
                 Y => SharedReg836_out);

   SharedReg837_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant15_0_impl_out,
                 Y => SharedReg837_out);

   SharedReg838_instance: Delay_34_DelayLength_22_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=22 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg837_out,
                 Y => SharedReg838_out);

   SharedReg839_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg838_out,
                 Y => SharedReg839_out);

   SharedReg840_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg839_out,
                 Y => SharedReg840_out);

   SharedReg841_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg840_out,
                 Y => SharedReg841_out);

   SharedReg842_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg841_out,
                 Y => SharedReg842_out);

   SharedReg843_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg842_out,
                 Y => SharedReg843_out);

   SharedReg844_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant7_0_impl_out,
                 Y => SharedReg844_out);

   SharedReg845_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg844_out,
                 Y => SharedReg845_out);

   SharedReg846_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant16_0_impl_out,
                 Y => SharedReg846_out);

   SharedReg847_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg846_out,
                 Y => SharedReg847_out);

   SharedReg848_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant8_0_impl_out,
                 Y => SharedReg848_out);

   SharedReg849_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg848_out,
                 Y => SharedReg849_out);

   SharedReg850_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg849_out,
                 Y => SharedReg850_out);

   SharedReg851_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg850_out,
                 Y => SharedReg851_out);

   SharedReg852_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg851_out,
                 Y => SharedReg852_out);

   SharedReg853_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant17_0_impl_out,
                 Y => SharedReg853_out);

   SharedReg854_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg853_out,
                 Y => SharedReg854_out);

   SharedReg855_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg854_out,
                 Y => SharedReg855_out);

   SharedReg856_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg855_out,
                 Y => SharedReg856_out);

   SharedReg857_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg856_out,
                 Y => SharedReg857_out);

   SharedReg858_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant9_0_impl_out,
                 Y => SharedReg858_out);

   SharedReg859_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg858_out,
                 Y => SharedReg859_out);

   SharedReg860_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant18_0_impl_out,
                 Y => SharedReg860_out);

   SharedReg861_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg860_out,
                 Y => SharedReg861_out);

   SharedReg862_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_0_impl_out,
                 Y => SharedReg862_out);

   SharedReg863_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_0_impl_out,
                 Y => SharedReg863_out);
end architecture;

