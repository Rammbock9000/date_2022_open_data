--------------------------------------------------------------------------------
--                         ModuloCounter_13_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_13_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of ModuloCounter_13_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(3 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 12 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2371584
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2371584 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2371584 is
signal XX_m2371585 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m2371585 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m2371585 <= X ;
   YY_m2371585 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_33_f500_uid2371588
--                   (IntAdderClassical_33_f500_uid2371590)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid2371588 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid2371588 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2371584 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid2371588 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid2371584  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
      RoundingAdder: IntAdder_33_f500_uid2371588  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_13_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_13_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_13_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
         iS_9 when "1001",
         iS_10 when "1010",
         iS_11 when "1011",
         iS_12 when "1100",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid2373455_RightShifter
--                (RightShifter_24_by_max_26_F250_uid2373457)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2373455_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2373455_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid2373460
--                  (IntAdderAlternative_27_f250_uid2373464)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid2373460 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid2373460 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid2373467
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid2373467 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid2373467 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid2373470
--                   (IntAdderClassical_34_f250_uid2373472)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid2373470 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid2373470 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid2373455
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2373455 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2373455 is
   component FPAdd_8_23_uid2373455_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid2373460 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid2373467 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid2373470 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid2373455_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid2373460  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid2373467  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid2373470  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid2373455 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid2373455  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_11_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_11_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_11_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
         iS_9 when "1001",
         iS_10 when "1010",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_12_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_12_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_12_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
         iS_9 when "1001",
         iS_10 when "1010",
         iS_11 when "1011",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid2374379_RightShifter
--                (RightShifter_24_by_max_26_F250_uid2374381)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2374379_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2374379_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid2374384
--                  (IntAdderAlternative_27_f250_uid2374388)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid2374384 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid2374384 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid2374391
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid2374391 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid2374391 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid2374394
--                   (IntAdderClassical_34_f250_uid2374396)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid2374394 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid2374394 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid2374379
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid2374379 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid2374379 is
   component FPAdd_8_23_uid2374379_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid2374384 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid2374391 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid2374394 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid2374379_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid2374384  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid2374391  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid2374394  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
   component FPAdd_8_23_uid2374379 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= (Y(Y'length-1 downto Y'length-2)) & (not Y(Y'length-3)) & Y(Y'length-4 downto 0);
   FPAddSubOp_instance: FPAdd_8_23_uid2374379  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_10_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_10_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(3 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_10_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "0000",
         iS_1 when "0001",
         iS_2 when "0010",
         iS_3 when "0011",
         iS_4 when "0100",
         iS_5 when "0101",
         iS_6 when "0110",
         iS_7 when "0111",
         iS_8 when "1000",
         iS_9 when "1001",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                      Constant_float_8_23_1_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111111100000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                            SelFunctionTable_r8
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
entity SelFunctionTable_r8 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(6 downto 0);
          Y : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of SelFunctionTable_r8 is
begin
  with X select  Y <= 
   "0000" when "0000000",
   "0000" when "0000001",
   "0000" when "0000010",
   "0000" when "0000011",
   "0001" when "0000100",
   "0001" when "0000101",
   "0001" when "0000110",
   "0001" when "0000111",
   "0001" when "0001000",
   "0001" when "0001001",
   "0001" when "0001010",
   "0001" when "0001011",
   "0010" when "0001100",
   "0010" when "0001101",
   "0010" when "0001110",
   "0010" when "0001111",
   "0011" when "0010000",
   "0011" when "0010001",
   "0010" when "0010010",
   "0010" when "0010011",
   "0011" when "0010100",
   "0011" when "0010101",
   "0011" when "0010110",
   "0011" when "0010111",
   "0100" when "0011000",
   "0100" when "0011001",
   "0011" when "0011010",
   "0011" when "0011011",
   "0101" when "0011100",
   "0100" when "0011101",
   "0100" when "0011110",
   "0100" when "0011111",
   "0101" when "0100000",
   "0101" when "0100001",
   "0101" when "0100010",
   "0100" when "0100011",
   "0110" when "0100100",
   "0110" when "0100101",
   "0101" when "0100110",
   "0101" when "0100111",
   "0111" when "0101000",
   "0110" when "0101001",
   "0110" when "0101010",
   "0101" when "0101011",
   "0111" when "0101100",
   "0111" when "0101101",
   "0110" when "0101110",
   "0110" when "0101111",
   "0111" when "0110000",
   "0111" when "0110001",
   "0111" when "0110010",
   "0110" when "0110011",
   "0111" when "0110100",
   "0111" when "0110101",
   "0111" when "0110110",
   "0111" when "0110111",
   "0111" when "0111000",
   "0111" when "0111001",
   "0111" when "0111010",
   "0111" when "0111011",
   "0111" when "0111100",
   "0111" when "0111101",
   "0111" when "0111110",
   "0111" when "0111111",
   "1001" when "1000000",
   "1001" when "1000001",
   "1001" when "1000010",
   "1001" when "1000011",
   "1001" when "1000100",
   "1001" when "1000101",
   "1001" when "1000110",
   "1001" when "1000111",
   "1001" when "1001000",
   "1001" when "1001001",
   "1001" when "1001010",
   "1001" when "1001011",
   "1001" when "1001100",
   "1001" when "1001101",
   "1001" when "1001110",
   "1001" when "1001111",
   "1001" when "1010000",
   "1001" when "1010001",
   "1010" when "1010010",
   "1010" when "1010011",
   "1001" when "1010100",
   "1010" when "1010101",
   "1010" when "1010110",
   "1010" when "1010111",
   "1010" when "1011000",
   "1010" when "1011001",
   "1011" when "1011010",
   "1011" when "1011011",
   "1011" when "1011100",
   "1011" when "1011101",
   "1011" when "1011110",
   "1011" when "1011111",
   "1011" when "1100000",
   "1011" when "1100001",
   "1100" when "1100010",
   "1100" when "1100011",
   "1100" when "1100100",
   "1100" when "1100101",
   "1100" when "1100110",
   "1100" when "1100111",
   "1100" when "1101000",
   "1101" when "1101001",
   "1101" when "1101010",
   "1101" when "1101011",
   "1101" when "1101100",
   "1101" when "1101101",
   "1101" when "1101110",
   "1101" when "1101111",
   "1110" when "1110000",
   "1110" when "1110001",
   "1110" when "1110010",
   "1110" when "1110011",
   "1110" when "1110100",
   "1110" when "1110101",
   "1110" when "1110110",
   "1110" when "1110111",
   "1111" when "1111000",
   "1111" when "1111001",
   "1111" when "1111010",
   "1111" when "1111011",
   "1111" when "1111100",
   "1111" when "1111101",
   "1111" when "1111110",
   "1111" when "1111111",
   "----" when others;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
   component SelFunctionTable_r8 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(6 downto 0);
             Y : out std_logic_vector(3 downto 0)   );
   end component;

signal partialFX : std_logic_vector(23 downto 0) := (others => '0');
signal partialFY : std_logic_vector(23 downto 0) := (others => '0');
signal expR0, expR0_d1, expR0_d2, expR0_d3, expR0_d4, expR0_d5, expR0_d6, expR0_d7, expR0_d8, expR0_d9, expR0_d10, expR0_d11 : std_logic_vector(9 downto 0) := (others => '0');
signal sR, sR_d1, sR_d2, sR_d3, sR_d4, sR_d5, sR_d6, sR_d7, sR_d8, sR_d9, sR_d10, sR_d11, sR_d12 : std_logic := '0';
signal exnXY : std_logic_vector(3 downto 0) := (others => '0');
signal exnR0, exnR0_d1, exnR0_d2, exnR0_d3, exnR0_d4, exnR0_d5, exnR0_d6, exnR0_d7, exnR0_d8, exnR0_d9, exnR0_d10, exnR0_d11, exnR0_d12 : std_logic_vector(1 downto 0) := (others => '0');
signal fY, fY_d1, fY_d2, fY_d3, fY_d4, fY_d5, fY_d6, fY_d7, fY_d8, fY_d9 : std_logic_vector(25 downto 0) := (others => '0');
signal fX : std_logic_vector(26 downto 0) := (others => '0');
signal w9, w9_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel9 : std_logic_vector(6 downto 0) := (others => '0');
signal q9, q9_d1, q9_d2, q9_d3, q9_d4, q9_d5, q9_d6, q9_d7, q9_d8, q9_d9 : std_logic_vector(3 downto 0) := (others => '0');
signal w9pad : std_logic_vector(29 downto 0) := (others => '0');
signal w8fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec8 : std_logic_vector(29 downto 0) := (others => '0');
signal w8full : std_logic_vector(29 downto 0) := (others => '0');
signal w8, w8_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel8 : std_logic_vector(6 downto 0) := (others => '0');
signal q8, q8_d1, q8_d2, q8_d3, q8_d4, q8_d5, q8_d6, q8_d7, q8_d8 : std_logic_vector(3 downto 0) := (others => '0');
signal w8pad : std_logic_vector(29 downto 0) := (others => '0');
signal w7fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec7 : std_logic_vector(29 downto 0) := (others => '0');
signal w7full : std_logic_vector(29 downto 0) := (others => '0');
signal w7, w7_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel7 : std_logic_vector(6 downto 0) := (others => '0');
signal q7, q7_d1, q7_d2, q7_d3, q7_d4, q7_d5, q7_d6, q7_d7 : std_logic_vector(3 downto 0) := (others => '0');
signal w7pad : std_logic_vector(29 downto 0) := (others => '0');
signal w6fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec6 : std_logic_vector(29 downto 0) := (others => '0');
signal w6full : std_logic_vector(29 downto 0) := (others => '0');
signal w6, w6_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel6 : std_logic_vector(6 downto 0) := (others => '0');
signal q6, q6_d1, q6_d2, q6_d3, q6_d4, q6_d5, q6_d6 : std_logic_vector(3 downto 0) := (others => '0');
signal w6pad : std_logic_vector(29 downto 0) := (others => '0');
signal w5fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec5 : std_logic_vector(29 downto 0) := (others => '0');
signal w5full : std_logic_vector(29 downto 0) := (others => '0');
signal w5, w5_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel5 : std_logic_vector(6 downto 0) := (others => '0');
signal q5, q5_d1, q5_d2, q5_d3, q5_d4, q5_d5 : std_logic_vector(3 downto 0) := (others => '0');
signal w5pad : std_logic_vector(29 downto 0) := (others => '0');
signal w4fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec4 : std_logic_vector(29 downto 0) := (others => '0');
signal w4full : std_logic_vector(29 downto 0) := (others => '0');
signal w4, w4_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel4 : std_logic_vector(6 downto 0) := (others => '0');
signal q4, q4_d1, q4_d2, q4_d3, q4_d4 : std_logic_vector(3 downto 0) := (others => '0');
signal w4pad : std_logic_vector(29 downto 0) := (others => '0');
signal w3fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec3 : std_logic_vector(29 downto 0) := (others => '0');
signal w3full : std_logic_vector(29 downto 0) := (others => '0');
signal w3, w3_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel3 : std_logic_vector(6 downto 0) := (others => '0');
signal q3, q3_d1, q3_d2, q3_d3 : std_logic_vector(3 downto 0) := (others => '0');
signal w3pad : std_logic_vector(29 downto 0) := (others => '0');
signal w2fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec2 : std_logic_vector(29 downto 0) := (others => '0');
signal w2full : std_logic_vector(29 downto 0) := (others => '0');
signal w2, w2_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel2 : std_logic_vector(6 downto 0) := (others => '0');
signal q2, q2_d1, q2_d2 : std_logic_vector(3 downto 0) := (others => '0');
signal w2pad : std_logic_vector(29 downto 0) := (others => '0');
signal w1fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec1 : std_logic_vector(29 downto 0) := (others => '0');
signal w1full : std_logic_vector(29 downto 0) := (others => '0');
signal w1, w1_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal sel1 : std_logic_vector(6 downto 0) := (others => '0');
signal q1, q1_d1 : std_logic_vector(3 downto 0) := (others => '0');
signal w1pad : std_logic_vector(29 downto 0) := (others => '0');
signal w0fulla : std_logic_vector(29 downto 0) := (others => '0');
signal fYdec0 : std_logic_vector(29 downto 0) := (others => '0');
signal w0full : std_logic_vector(29 downto 0) := (others => '0');
signal w0, w0_d1 : std_logic_vector(28 downto 0) := (others => '0');
signal q0 : std_logic_vector(3 downto 0) := (others => '0');
signal qP9 : std_logic_vector(2 downto 0) := (others => '0');
signal qM9 : std_logic_vector(2 downto 0) := (others => '0');
signal qP8 : std_logic_vector(2 downto 0) := (others => '0');
signal qM8 : std_logic_vector(2 downto 0) := (others => '0');
signal qP7 : std_logic_vector(2 downto 0) := (others => '0');
signal qM7 : std_logic_vector(2 downto 0) := (others => '0');
signal qP6 : std_logic_vector(2 downto 0) := (others => '0');
signal qM6 : std_logic_vector(2 downto 0) := (others => '0');
signal qP5 : std_logic_vector(2 downto 0) := (others => '0');
signal qM5 : std_logic_vector(2 downto 0) := (others => '0');
signal qP4 : std_logic_vector(2 downto 0) := (others => '0');
signal qM4 : std_logic_vector(2 downto 0) := (others => '0');
signal qP3 : std_logic_vector(2 downto 0) := (others => '0');
signal qM3 : std_logic_vector(2 downto 0) := (others => '0');
signal qP2 : std_logic_vector(2 downto 0) := (others => '0');
signal qM2 : std_logic_vector(2 downto 0) := (others => '0');
signal qP1 : std_logic_vector(2 downto 0) := (others => '0');
signal qM1 : std_logic_vector(2 downto 0) := (others => '0');
signal qP0 : std_logic_vector(2 downto 0) := (others => '0');
signal qM0 : std_logic_vector(2 downto 0) := (others => '0');
signal qP : std_logic_vector(29 downto 0) := (others => '0');
signal qM : std_logic_vector(29 downto 0) := (others => '0');
signal fR0, fR0_d1 : std_logic_vector(29 downto 0) := (others => '0');
signal fR : std_logic_vector(28 downto 0) := (others => '0');
signal fRn1, fRn1_d1 : std_logic_vector(26 downto 0) := (others => '0');
signal expR1, expR1_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal round, round_d1 : std_logic := '0';
signal expfrac : std_logic_vector(32 downto 0) := (others => '0');
signal expfracR : std_logic_vector(32 downto 0) := (others => '0');
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
signal exnRfinal : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            expR0_d1 <=  expR0;
            expR0_d2 <=  expR0_d1;
            expR0_d3 <=  expR0_d2;
            expR0_d4 <=  expR0_d3;
            expR0_d5 <=  expR0_d4;
            expR0_d6 <=  expR0_d5;
            expR0_d7 <=  expR0_d6;
            expR0_d8 <=  expR0_d7;
            expR0_d9 <=  expR0_d8;
            expR0_d10 <=  expR0_d9;
            expR0_d11 <=  expR0_d10;
            sR_d1 <=  sR;
            sR_d2 <=  sR_d1;
            sR_d3 <=  sR_d2;
            sR_d4 <=  sR_d3;
            sR_d5 <=  sR_d4;
            sR_d6 <=  sR_d5;
            sR_d7 <=  sR_d6;
            sR_d8 <=  sR_d7;
            sR_d9 <=  sR_d8;
            sR_d10 <=  sR_d9;
            sR_d11 <=  sR_d10;
            sR_d12 <=  sR_d11;
            exnR0_d1 <=  exnR0;
            exnR0_d2 <=  exnR0_d1;
            exnR0_d3 <=  exnR0_d2;
            exnR0_d4 <=  exnR0_d3;
            exnR0_d5 <=  exnR0_d4;
            exnR0_d6 <=  exnR0_d5;
            exnR0_d7 <=  exnR0_d6;
            exnR0_d8 <=  exnR0_d7;
            exnR0_d9 <=  exnR0_d8;
            exnR0_d10 <=  exnR0_d9;
            exnR0_d11 <=  exnR0_d10;
            exnR0_d12 <=  exnR0_d11;
            fY_d1 <=  fY;
            fY_d2 <=  fY_d1;
            fY_d3 <=  fY_d2;
            fY_d4 <=  fY_d3;
            fY_d5 <=  fY_d4;
            fY_d6 <=  fY_d5;
            fY_d7 <=  fY_d6;
            fY_d8 <=  fY_d7;
            fY_d9 <=  fY_d8;
            w9_d1 <=  w9;
            q9_d1 <=  q9;
            q9_d2 <=  q9_d1;
            q9_d3 <=  q9_d2;
            q9_d4 <=  q9_d3;
            q9_d5 <=  q9_d4;
            q9_d6 <=  q9_d5;
            q9_d7 <=  q9_d6;
            q9_d8 <=  q9_d7;
            q9_d9 <=  q9_d8;
            w8_d1 <=  w8;
            q8_d1 <=  q8;
            q8_d2 <=  q8_d1;
            q8_d3 <=  q8_d2;
            q8_d4 <=  q8_d3;
            q8_d5 <=  q8_d4;
            q8_d6 <=  q8_d5;
            q8_d7 <=  q8_d6;
            q8_d8 <=  q8_d7;
            w7_d1 <=  w7;
            q7_d1 <=  q7;
            q7_d2 <=  q7_d1;
            q7_d3 <=  q7_d2;
            q7_d4 <=  q7_d3;
            q7_d5 <=  q7_d4;
            q7_d6 <=  q7_d5;
            q7_d7 <=  q7_d6;
            w6_d1 <=  w6;
            q6_d1 <=  q6;
            q6_d2 <=  q6_d1;
            q6_d3 <=  q6_d2;
            q6_d4 <=  q6_d3;
            q6_d5 <=  q6_d4;
            q6_d6 <=  q6_d5;
            w5_d1 <=  w5;
            q5_d1 <=  q5;
            q5_d2 <=  q5_d1;
            q5_d3 <=  q5_d2;
            q5_d4 <=  q5_d3;
            q5_d5 <=  q5_d4;
            w4_d1 <=  w4;
            q4_d1 <=  q4;
            q4_d2 <=  q4_d1;
            q4_d3 <=  q4_d2;
            q4_d4 <=  q4_d3;
            w3_d1 <=  w3;
            q3_d1 <=  q3;
            q3_d2 <=  q3_d1;
            q3_d3 <=  q3_d2;
            w2_d1 <=  w2;
            q2_d1 <=  q2;
            q2_d2 <=  q2_d1;
            w1_d1 <=  w1;
            q1_d1 <=  q1;
            w0_d1 <=  w0;
            fR0_d1 <=  fR0;
            fRn1_d1 <=  fRn1;
            expR1_d1 <=  expR1;
            round_d1 <=  round;
         end if;
      end process;
   partialFX <= "1" & X(22 downto 0);
   partialFY <= "1" & Y(22 downto 0);
   -- exponent difference, sign and exception combination computed early, to have less bits to pipeline
   expR0 <= ("00" & X(30 downto 23)) - ("00" & Y(30 downto 23));
   sR <= X(31) xor Y(31);
   -- early exception handling 
   exnXY <= X(33 downto 32) & Y(33 downto 32);
   with exnXY select
      exnR0 <= 
         "01"  when "0101",                   -- normal
         "00"  when "0001" | "0010" | "0110", -- zero
         "10"  when "0100" | "1000" | "1001", -- overflow
         "11"  when others;                   -- NaN
    -- Prescaling
   with partialFY (22 downto 21) select
      fY <= 
         ("0" & partialFY & "0") + (partialFY & "00") when "00",
         ("00" & partialFY) + (partialFY & "00") when "01",
         partialFY &"00" when others;
   with partialFY (22 downto 21) select
      fX <= 
         ("00" & partialFX & "0") + ("0" & partialFX & "00") when "00",
         ("000" & partialFX) + ("0" & partialFX & "00") when "01",
         "0" & partialFX &"00" when others;
   w9 <=  "00" & fX;
   ----------------Synchro barrier, entering cycle 1----------------
   sel9 <= w9_d1(28 downto 24) & fY_d1(23 downto 22);
   SelFunctionTable9: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel9,
                 Y => q9);
   w9pad <= w9_d1 & '0';
   with q9(1 downto 0) select 
   w8fulla <= 
      w9pad - ("0000" & fY_d1)			when "01",
      w9pad + ("0000" & fY_d1)			when "11",
      w9pad + ("000" & fY_d1 & "0")	  when "10",
      w9pad 			   		  when others;
   with q9(3 downto 1) select 
   fYdec8 <= 
      ("00" & fY_d1 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d1 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q9(3) select
   w8full <= 
      w8fulla - fYdec8			when '0',
      w8fulla + fYdec8			when others;
   w8 <= w8full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 2----------------
   sel8 <= w8_d1(28 downto 24) & fY_d2(23 downto 22);
   SelFunctionTable8: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel8,
                 Y => q8);
   w8pad <= w8_d1 & '0';
   with q8(1 downto 0) select 
   w7fulla <= 
      w8pad - ("0000" & fY_d2)			when "01",
      w8pad + ("0000" & fY_d2)			when "11",
      w8pad + ("000" & fY_d2 & "0")	  when "10",
      w8pad 			   		  when others;
   with q8(3 downto 1) select 
   fYdec7 <= 
      ("00" & fY_d2 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d2 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q8(3) select
   w7full <= 
      w7fulla - fYdec7			when '0',
      w7fulla + fYdec7			when others;
   w7 <= w7full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 3----------------
   sel7 <= w7_d1(28 downto 24) & fY_d3(23 downto 22);
   SelFunctionTable7: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel7,
                 Y => q7);
   w7pad <= w7_d1 & '0';
   with q7(1 downto 0) select 
   w6fulla <= 
      w7pad - ("0000" & fY_d3)			when "01",
      w7pad + ("0000" & fY_d3)			when "11",
      w7pad + ("000" & fY_d3 & "0")	  when "10",
      w7pad 			   		  when others;
   with q7(3 downto 1) select 
   fYdec6 <= 
      ("00" & fY_d3 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d3 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q7(3) select
   w6full <= 
      w6fulla - fYdec6			when '0',
      w6fulla + fYdec6			when others;
   w6 <= w6full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 4----------------
   sel6 <= w6_d1(28 downto 24) & fY_d4(23 downto 22);
   SelFunctionTable6: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel6,
                 Y => q6);
   w6pad <= w6_d1 & '0';
   with q6(1 downto 0) select 
   w5fulla <= 
      w6pad - ("0000" & fY_d4)			when "01",
      w6pad + ("0000" & fY_d4)			when "11",
      w6pad + ("000" & fY_d4 & "0")	  when "10",
      w6pad 			   		  when others;
   with q6(3 downto 1) select 
   fYdec5 <= 
      ("00" & fY_d4 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d4 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q6(3) select
   w5full <= 
      w5fulla - fYdec5			when '0',
      w5fulla + fYdec5			when others;
   w5 <= w5full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 5----------------
   sel5 <= w5_d1(28 downto 24) & fY_d5(23 downto 22);
   SelFunctionTable5: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel5,
                 Y => q5);
   w5pad <= w5_d1 & '0';
   with q5(1 downto 0) select 
   w4fulla <= 
      w5pad - ("0000" & fY_d5)			when "01",
      w5pad + ("0000" & fY_d5)			when "11",
      w5pad + ("000" & fY_d5 & "0")	  when "10",
      w5pad 			   		  when others;
   with q5(3 downto 1) select 
   fYdec4 <= 
      ("00" & fY_d5 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d5 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q5(3) select
   w4full <= 
      w4fulla - fYdec4			when '0',
      w4fulla + fYdec4			when others;
   w4 <= w4full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 6----------------
   sel4 <= w4_d1(28 downto 24) & fY_d6(23 downto 22);
   SelFunctionTable4: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel4,
                 Y => q4);
   w4pad <= w4_d1 & '0';
   with q4(1 downto 0) select 
   w3fulla <= 
      w4pad - ("0000" & fY_d6)			when "01",
      w4pad + ("0000" & fY_d6)			when "11",
      w4pad + ("000" & fY_d6 & "0")	  when "10",
      w4pad 			   		  when others;
   with q4(3 downto 1) select 
   fYdec3 <= 
      ("00" & fY_d6 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d6 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q4(3) select
   w3full <= 
      w3fulla - fYdec3			when '0',
      w3fulla + fYdec3			when others;
   w3 <= w3full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 7----------------
   sel3 <= w3_d1(28 downto 24) & fY_d7(23 downto 22);
   SelFunctionTable3: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel3,
                 Y => q3);
   w3pad <= w3_d1 & '0';
   with q3(1 downto 0) select 
   w2fulla <= 
      w3pad - ("0000" & fY_d7)			when "01",
      w3pad + ("0000" & fY_d7)			when "11",
      w3pad + ("000" & fY_d7 & "0")	  when "10",
      w3pad 			   		  when others;
   with q3(3 downto 1) select 
   fYdec2 <= 
      ("00" & fY_d7 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d7 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q3(3) select
   w2full <= 
      w2fulla - fYdec2			when '0',
      w2fulla + fYdec2			when others;
   w2 <= w2full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 8----------------
   sel2 <= w2_d1(28 downto 24) & fY_d8(23 downto 22);
   SelFunctionTable2: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel2,
                 Y => q2);
   w2pad <= w2_d1 & '0';
   with q2(1 downto 0) select 
   w1fulla <= 
      w2pad - ("0000" & fY_d8)			when "01",
      w2pad + ("0000" & fY_d8)			when "11",
      w2pad + ("000" & fY_d8 & "0")	  when "10",
      w2pad 			   		  when others;
   with q2(3 downto 1) select 
   fYdec1 <= 
      ("00" & fY_d8 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d8 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q2(3) select
   w1full <= 
      w1fulla - fYdec1			when '0',
      w1fulla + fYdec1			when others;
   w1 <= w1full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 9----------------
   sel1 <= w1_d1(28 downto 24) & fY_d9(23 downto 22);
   SelFunctionTable1: SelFunctionTable_r8  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => sel1,
                 Y => q1);
   w1pad <= w1_d1 & '0';
   with q1(1 downto 0) select 
   w0fulla <= 
      w1pad - ("0000" & fY_d9)			when "01",
      w1pad + ("0000" & fY_d9)			when "11",
      w1pad + ("000" & fY_d9 & "0")	  when "10",
      w1pad 			   		  when others;
   with q1(3 downto 1) select 
   fYdec0 <= 
      ("00" & fY_d9 & "00")			when "001" | "010" | "110"| "101",
      ("0" & fY_d9 & "000")			when "011"| "100",
      (29 downto 0 => '0')when others;
   with q1(3) select
   w0full <= 
      w0fulla - fYdec0			when '0',
      w0fulla + fYdec0			when others;
   w0 <= w0full(26 downto 0) & "00";
   ----------------Synchro barrier, entering cycle 10----------------
   q0(3 downto 0) <= "0000" when  w0_d1 = (28 downto 0 => '0')
                else w0_d1(28) & "010";
   qP9 <=      q9_d9(2 downto 0);
   qM9 <=      q9_d9(3) & "00";
   qP8 <=      q8_d8(2 downto 0);
   qM8 <=      q8_d8(3) & "00";
   qP7 <=      q7_d7(2 downto 0);
   qM7 <=      q7_d7(3) & "00";
   qP6 <=      q6_d6(2 downto 0);
   qM6 <=      q6_d6(3) & "00";
   qP5 <=      q5_d5(2 downto 0);
   qM5 <=      q5_d5(3) & "00";
   qP4 <=      q4_d4(2 downto 0);
   qM4 <=      q4_d4(3) & "00";
   qP3 <=      q3_d3(2 downto 0);
   qM3 <=      q3_d3(3) & "00";
   qP2 <=      q2_d2(2 downto 0);
   qM2 <=      q2_d2(3) & "00";
   qP1 <=      q1_d1(2 downto 0);
   qM1 <=      q1_d1(3) & "00";
   qP0 <= q0(2 downto 0);
   qM0 <= q0(3)  & "00";
   qP <= qP9 & qP8 & qP7 & qP6 & qP5 & qP4 & qP3 & qP2 & qP1 & qP0;
   qM <= qM9(1 downto 0) & qM8 & qM7 & qM6 & qM5 & qM4 & qM3 & qM2 & qM1 & qM0 & "0";
   fR0 <= qP - qM;
   ----------------Synchro barrier, entering cycle 11----------------
   fR <= fR0_d1(29 downto 2) & (fR0_d1(0) or fR0_d1(1)); 
   -- normalisation
   with fR(27) select
      fRn1 <= fR(27 downto 2) & (fR(0) or fR(1)) when '1',
              fR(26 downto 0)          when others;
   expR1 <= expR0_d11 + ("000" & (6 downto 1 => '1') & fR(27)); -- add back bias
   round <= fRn1(2) and (fRn1(0) or fRn1(1) or fRn1(3)); -- fRn1(0) is the sticky bit
   ----------------Synchro barrier, entering cycle 12----------------
   -- final rounding
   expfrac <= expR1_d1 & fRn1_d1(25 downto 3) ;
   expfracR <= expfrac + ((32 downto 1 => '0') & round_d1);
   exnR <=      "00"  when expfracR(32) = '1'   -- underflow
           else "10"  when  expfracR(32 downto 31) =  "01" -- overflow
           else "01";      -- 00, normal case
   with exnR0_d12 select
      exnRfinal <= 
         exnR   when "01", -- normal
         exnR0_d12  when others;
   R <= exnRfinal & sR_d12 & expfracR(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_6_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_6_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(2 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_6_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000",
         iS_1 when "001",
         iS_2 when "010",
         iS_3 when "011",
         iS_4 when "100",
         iS_5 when "101",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_348_mult_8en9_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_348_mult_8en9_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_348_mult_8en9_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100110110001110101101010011000001";
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      Y <= s7;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 56 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      Y <= s55;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 24 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      Y <= s23;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 50 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      Y <= s49;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 19 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      Y <= s18;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      Y <= s13;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      Y <= s8;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      Y <= s11;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 39 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      Y <= s38;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 18 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      Y <= s17;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 27 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      Y <= s26;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 42 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      Y <= s41;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_95_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 95 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_95_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_95_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      Y <= s94;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_87_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 87 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_87_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_87_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      Y <= s86;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_85_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 85 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_85_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_85_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      Y <= s84;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_97_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 97 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_97_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_97_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      Y <= s96;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 49 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      Y <= s48;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 64 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      Y <= s63;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      Y <= s10;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 65 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      Y <= s64;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_68_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 68 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_68_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_68_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      Y <= s67;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 15 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      Y <= s14;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 45 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      Y <= s44;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 29 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      Y <= s28;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      Y <= s9;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 35 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      Y <= s34;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 57 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      Y <= s56;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      Y <= s12;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 61 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      Y <= s60;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 40 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      Y <= s39;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 36 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      Y <= s35;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 43 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      Y <= s42;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 44 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      Y <= s43;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Add141_5_impl_0_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add141_5_impl_0_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add141_5_impl_0_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0110" when "0000",
      "1000" when "0001",
      "0011" when "0010",
      "0000" when "0011",
      "1001" when "0100",
      "0001" when "0101",
      "0101" when "0110",
      "1010" when "0111",
      "0000" when "1000",
      "0000" when "1001",
      "0010" when "1010",
      "0100" when "1011",
      "0111" when "1100",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Add141_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add141_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add141_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Add141_5_impl_0_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Add141_5_impl_0_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Add141_5_impl_1_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add141_5_impl_1_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add141_5_impl_1_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0010" when "0000",
      "1000" when "0001",
      "0101" when "0010",
      "1010" when "0011",
      "0111" when "0100",
      "0011" when "0101",
      "0001" when "0110",
      "1001" when "0111",
      "0000" when "1000",
      "0000" when "1001",
      "0100" when "1010",
      "0000" when "1011",
      "0110" when "1100",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Add141_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add141_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add141_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Add141_5_impl_1_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Add141_5_impl_1_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product62_5_impl_0_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product62_5_impl_0_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product62_5_impl_0_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "1001" when "0000",
      "0000" when "0001",
      "0100" when "0010",
      "1011" when "0011",
      "1010" when "0100",
      "0111" when "0101",
      "0010" when "0110",
      "0101" when "0111",
      "1000" when "1000",
      "0110" when "1001",
      "0001" when "1010",
      "0000" when "1011",
      "0011" when "1100",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product62_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product62_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product62_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product62_5_impl_0_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product62_5_impl_0_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product62_5_impl_1_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product62_5_impl_1_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product62_5_impl_1_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0101" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0110" when "0011",
      "0100" when "0100",
      "1010" when "0101",
      "0001" when "0110",
      "1000" when "0111",
      "0111" when "1000",
      "1001" when "1001",
      "0011" when "1010",
      "0010" when "1011",
      "1011" when "1100",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product62_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product62_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product62_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product62_5_impl_1_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product62_5_impl_1_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add10_5_impl_0_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add10_5_impl_0_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add10_5_impl_0_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0101" when "0000",
      "0000" when "0001",
      "0010" when "0010",
      "0000" when "0011",
      "1000" when "0100",
      "0100" when "0101",
      "0111" when "0110",
      "0001" when "0111",
      "0000" when "1000",
      "0000" when "1001",
      "0011" when "1010",
      "0110" when "1011",
      "1001" when "1100",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add10_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add10_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add10_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Add10_5_impl_0_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Add10_5_impl_0_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--           GenericLut_LUTData_MUX_Add10_5_impl_1_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add10_5_impl_1_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add10_5_impl_1_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "1000" when "0000",
      "0000" when "0001",
      "0001" when "0010",
      "1001" when "0011",
      "0000" when "0100",
      "0110" when "0101",
      "0100" when "0110",
      "0010" when "0111",
      "0000" when "1000",
      "0000" when "1001",
      "0111" when "1010",
      "0101" when "1011",
      "0011" when "1100",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--  GenericLut_LUTData_MUX_Add10_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Add10_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Add10_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Add10_5_impl_1_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Add10_5_impl_1_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "101" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "001" when "0101",
      "000" when "0110",
      "010" when "0111",
      "000" when "1000",
      "011" when "1001",
      "000" when "1010",
      "100" when "1011",
      "000" when "1100",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "000" when "0000",
      "101" when "0001",
      "000" when "0010",
      "000" when "0011",
      "000" when "0100",
      "001" when "0101",
      "000" when "0110",
      "010" when "0111",
      "000" when "1000",
      "011" when "1001",
      "000" when "1010",
      "100" when "1011",
      "000" when "1100",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product213_5_impl_0_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product213_5_impl_0_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product213_5_impl_0_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0000" when "0000",
      "0000" when "0001",
      "0011" when "0010",
      "1000" when "0011",
      "0111" when "0100",
      "0101" when "0101",
      "0100" when "0110",
      "0000" when "0111",
      "1001" when "1000",
      "0010" when "1001",
      "0000" when "1010",
      "0110" when "1011",
      "0001" when "1100",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product213_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product213_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product213_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product213_5_impl_0_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product213_5_impl_0_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--        GenericLut_LUTData_MUX_Product213_5_impl_1_LUT_wIn_4_wOut_4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product213_5_impl_1_LUT_wIn_4_wOut_4 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product213_5_impl_1_LUT_wIn_4_wOut_4 is
signal t_in : std_logic_vector(3 downto 0) := (others => '0');
signal t_out : std_logic_vector(3 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   with t_in select t_out <= 
      "0000" when "0000",
      "0000" when "0001",
      "1000" when "0010",
      "0101" when "0011",
      "0011" when "0100",
      "0110" when "0101",
      "0100" when "0110",
      "0000" when "0111",
      "0001" when "1000",
      "0111" when "1001",
      "0000" when "1010",
      "0010" when "1011",
      "1001" when "1100",
      "0000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product213_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product213_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(3 downto 0);
          Output : out std_logic_vector(3 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product213_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
   component GenericLut_LUTData_MUX_Product213_5_impl_1_LUT_wIn_4_wOut_4 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
   instLUT: GenericLut_LUTData_MUX_Product213_5_impl_1_LUT_wIn_4_wOut_4
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 28 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      Y <= s27;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 48 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      Y <= s47;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_78_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 78 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_78_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_78_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      Y <= s77;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 67 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      Y <= s66;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 38 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      Y <= s37;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 55 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      Y <= s54;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 53 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      Y <= s52;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 47 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      Y <= s46;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 63 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      Y <= s62;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 58 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      Y <= s57;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 62 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      Y <= s61;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_51_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 51 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_51_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_51_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      Y <= s50;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 52 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      Y <= s51;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 46 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      Y <= s45;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 17 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      Y <= s16;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 32 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      Y <= s31;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 30 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      Y <= s29;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 31 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      Y <= s30;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 26 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      Y <= s25;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_103_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 103 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_103_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_103_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      Y <= s102;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      Y <= s20;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          Ldiff_UU_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_UU_del_1_1 : in std_logic_vector(31 downto 0);
          Ldiff_UU_del_1_2 : in std_logic_vector(31 downto 0);
          Ldiff_UU_del_1_3 : in std_logic_vector(31 downto 0);
          Ldiff_UU_del_1_4 : in std_logic_vector(31 downto 0);
          Ldiff_UU_del_1_5 : in std_logic_vector(31 downto 0);
          Ldiff_UV_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_UV_del_1_1 : in std_logic_vector(31 downto 0);
          Ldiff_UV_del_1_2 : in std_logic_vector(31 downto 0);
          Ldiff_UV_del_1_3 : in std_logic_vector(31 downto 0);
          Ldiff_UV_del_1_4 : in std_logic_vector(31 downto 0);
          Ldiff_UV_del_1_5 : in std_logic_vector(31 downto 0);
          Ldiff_UW_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_UW_del_1_1 : in std_logic_vector(31 downto 0);
          Ldiff_UW_del_1_2 : in std_logic_vector(31 downto 0);
          Ldiff_UW_del_1_3 : in std_logic_vector(31 downto 0);
          Ldiff_UW_del_1_4 : in std_logic_vector(31 downto 0);
          Ldiff_UW_del_1_5 : in std_logic_vector(31 downto 0);
          Ldiff_VU_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_VU_del_1_1 : in std_logic_vector(31 downto 0);
          Ldiff_VU_del_1_2 : in std_logic_vector(31 downto 0);
          Ldiff_VU_del_1_3 : in std_logic_vector(31 downto 0);
          Ldiff_VU_del_1_4 : in std_logic_vector(31 downto 0);
          Ldiff_VU_del_1_5 : in std_logic_vector(31 downto 0);
          Ldiff_VV_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_VV_del_1_1 : in std_logic_vector(31 downto 0);
          Ldiff_VV_del_1_2 : in std_logic_vector(31 downto 0);
          Ldiff_VV_del_1_3 : in std_logic_vector(31 downto 0);
          Ldiff_VV_del_1_4 : in std_logic_vector(31 downto 0);
          Ldiff_VV_del_1_5 : in std_logic_vector(31 downto 0);
          Ldiff_VW_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_VW_del_1_1 : in std_logic_vector(31 downto 0);
          Ldiff_VW_del_1_2 : in std_logic_vector(31 downto 0);
          Ldiff_VW_del_1_3 : in std_logic_vector(31 downto 0);
          Ldiff_VW_del_1_4 : in std_logic_vector(31 downto 0);
          Ldiff_VW_del_1_5 : in std_logic_vector(31 downto 0);
          Ldiff_WU_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_WU_del_1_1 : in std_logic_vector(31 downto 0);
          Ldiff_WU_del_1_2 : in std_logic_vector(31 downto 0);
          Ldiff_WU_del_1_3 : in std_logic_vector(31 downto 0);
          Ldiff_WU_del_1_4 : in std_logic_vector(31 downto 0);
          Ldiff_WU_del_1_5 : in std_logic_vector(31 downto 0);
          Ldiff_WV_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_WV_del_1_1 : in std_logic_vector(31 downto 0);
          Ldiff_WV_del_1_2 : in std_logic_vector(31 downto 0);
          Ldiff_WV_del_1_3 : in std_logic_vector(31 downto 0);
          Ldiff_WV_del_1_4 : in std_logic_vector(31 downto 0);
          Ldiff_WV_del_1_5 : in std_logic_vector(31 downto 0);
          Ldiff_WW_del_1_0 : in std_logic_vector(31 downto 0);
          Ldiff_WW_del_1_1 : in std_logic_vector(31 downto 0);
          Ldiff_WW_del_1_2 : in std_logic_vector(31 downto 0);
          Ldiff_WW_del_1_3 : in std_logic_vector(31 downto 0);
          Ldiff_WW_del_1_4 : in std_logic_vector(31 downto 0);
          Ldiff_WW_del_1_5 : in std_logic_vector(31 downto 0);
          R_U_0 : in std_logic_vector(31 downto 0);
          R_U_1 : in std_logic_vector(31 downto 0);
          R_U_2 : in std_logic_vector(31 downto 0);
          R_U_3 : in std_logic_vector(31 downto 0);
          R_U_4 : in std_logic_vector(31 downto 0);
          R_U_5 : in std_logic_vector(31 downto 0);
          R_V_0 : in std_logic_vector(31 downto 0);
          R_V_1 : in std_logic_vector(31 downto 0);
          R_V_2 : in std_logic_vector(31 downto 0);
          R_V_3 : in std_logic_vector(31 downto 0);
          R_V_4 : in std_logic_vector(31 downto 0);
          R_V_5 : in std_logic_vector(31 downto 0);
          R_W_0 : in std_logic_vector(31 downto 0);
          R_W_1 : in std_logic_vector(31 downto 0);
          R_W_2 : in std_logic_vector(31 downto 0);
          R_W_3 : in std_logic_vector(31 downto 0);
          R_W_4 : in std_logic_vector(31 downto 0);
          R_W_5 : in std_logic_vector(31 downto 0);
          Inv_11_0 : out std_logic_vector(31 downto 0);
          Inv_11_1 : out std_logic_vector(31 downto 0);
          Inv_11_2 : out std_logic_vector(31 downto 0);
          Inv_11_3 : out std_logic_vector(31 downto 0);
          Inv_11_4 : out std_logic_vector(31 downto 0);
          Inv_11_5 : out std_logic_vector(31 downto 0);
          Inv_12_0 : out std_logic_vector(31 downto 0);
          Inv_12_1 : out std_logic_vector(31 downto 0);
          Inv_12_2 : out std_logic_vector(31 downto 0);
          Inv_12_3 : out std_logic_vector(31 downto 0);
          Inv_12_4 : out std_logic_vector(31 downto 0);
          Inv_12_5 : out std_logic_vector(31 downto 0);
          Inv_13_0 : out std_logic_vector(31 downto 0);
          Inv_13_1 : out std_logic_vector(31 downto 0);
          Inv_13_2 : out std_logic_vector(31 downto 0);
          Inv_13_3 : out std_logic_vector(31 downto 0);
          Inv_13_4 : out std_logic_vector(31 downto 0);
          Inv_13_5 : out std_logic_vector(31 downto 0);
          Inv_21_0 : out std_logic_vector(31 downto 0);
          Inv_21_1 : out std_logic_vector(31 downto 0);
          Inv_21_2 : out std_logic_vector(31 downto 0);
          Inv_21_3 : out std_logic_vector(31 downto 0);
          Inv_21_4 : out std_logic_vector(31 downto 0);
          Inv_21_5 : out std_logic_vector(31 downto 0);
          Inv_22_0 : out std_logic_vector(31 downto 0);
          Inv_22_1 : out std_logic_vector(31 downto 0);
          Inv_22_2 : out std_logic_vector(31 downto 0);
          Inv_22_3 : out std_logic_vector(31 downto 0);
          Inv_22_4 : out std_logic_vector(31 downto 0);
          Inv_22_5 : out std_logic_vector(31 downto 0);
          Inv_23_0 : out std_logic_vector(31 downto 0);
          Inv_23_1 : out std_logic_vector(31 downto 0);
          Inv_23_2 : out std_logic_vector(31 downto 0);
          Inv_23_3 : out std_logic_vector(31 downto 0);
          Inv_23_4 : out std_logic_vector(31 downto 0);
          Inv_23_5 : out std_logic_vector(31 downto 0);
          Inv_31_0 : out std_logic_vector(31 downto 0);
          Inv_31_1 : out std_logic_vector(31 downto 0);
          Inv_31_2 : out std_logic_vector(31 downto 0);
          Inv_31_3 : out std_logic_vector(31 downto 0);
          Inv_31_4 : out std_logic_vector(31 downto 0);
          Inv_31_5 : out std_logic_vector(31 downto 0);
          Inv_32_0 : out std_logic_vector(31 downto 0);
          Inv_32_1 : out std_logic_vector(31 downto 0);
          Inv_32_2 : out std_logic_vector(31 downto 0);
          Inv_32_3 : out std_logic_vector(31 downto 0);
          Inv_32_4 : out std_logic_vector(31 downto 0);
          Inv_32_5 : out std_logic_vector(31 downto 0);
          Inv_33_0 : out std_logic_vector(31 downto 0);
          Inv_33_1 : out std_logic_vector(31 downto 0);
          Inv_33_2 : out std_logic_vector(31 downto 0);
          Inv_33_3 : out std_logic_vector(31 downto 0);
          Inv_33_4 : out std_logic_vector(31 downto 0);
          Inv_33_5 : out std_logic_vector(31 downto 0);
          Inv_41_0 : out std_logic_vector(31 downto 0);
          Inv_41_1 : out std_logic_vector(31 downto 0);
          Inv_41_2 : out std_logic_vector(31 downto 0);
          Inv_41_3 : out std_logic_vector(31 downto 0);
          Inv_41_4 : out std_logic_vector(31 downto 0);
          Inv_41_5 : out std_logic_vector(31 downto 0);
          Inv_42_0 : out std_logic_vector(31 downto 0);
          Inv_42_1 : out std_logic_vector(31 downto 0);
          Inv_42_2 : out std_logic_vector(31 downto 0);
          Inv_42_3 : out std_logic_vector(31 downto 0);
          Inv_42_4 : out std_logic_vector(31 downto 0);
          Inv_42_5 : out std_logic_vector(31 downto 0);
          Inv_43_0 : out std_logic_vector(31 downto 0);
          Inv_43_1 : out std_logic_vector(31 downto 0);
          Inv_43_2 : out std_logic_vector(31 downto 0);
          Inv_43_3 : out std_logic_vector(31 downto 0);
          Inv_43_4 : out std_logic_vector(31 downto 0);
          Inv_43_5 : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_13_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(3 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_13_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_11_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_12_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_10_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(3 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Constant_float_8_23_1_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_6_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(2 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Constant_float_8_23_348_mult_8en9_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_95_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_87_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_85_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_97_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_68_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add141_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add141_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product62_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product62_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add10_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Add10_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product213_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product213_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(3 downto 0);
             Output : out std_logic_vector(3 downto 0)   );
   end component;

   component Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_78_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_51_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_103_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount131_out : std_logic_vector(3 downto 0) := (others => '0');
signal Ldiff_UU_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UU_del_1_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UU_del_1_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UU_del_1_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UU_del_1_4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UU_del_1_5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UV_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UV_del_1_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UV_del_1_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UV_del_1_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UV_del_1_4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UV_del_1_5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UW_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UW_del_1_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UW_del_1_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UW_del_1_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UW_del_1_4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UW_del_1_5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VU_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VU_del_1_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VU_del_1_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VU_del_1_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VU_del_1_4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VU_del_1_5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VV_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VV_del_1_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VV_del_1_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VV_del_1_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VV_del_1_4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VV_del_1_5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VW_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VW_del_1_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VW_del_1_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VW_del_1_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VW_del_1_4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_VW_del_1_5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WU_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WU_del_1_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WU_del_1_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WU_del_1_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WU_del_1_4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WU_del_1_5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WV_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WV_del_1_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WV_del_1_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WV_del_1_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WV_del_1_4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WV_del_1_5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WW_del_1_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WW_del_1_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WW_del_1_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WW_del_1_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WW_del_1_4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_WW_del_1_5_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_U_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_U_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_U_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_U_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_U_4_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_U_5_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_V_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_V_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_V_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_V_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_V_4_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_V_5_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_W_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_W_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_W_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_W_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_W_4_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_W_5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product108_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product108_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product110_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product110_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product109_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product109_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product109_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product109_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product109_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product109_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product109_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product111_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product111_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product210_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product210_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product310_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product310_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product410_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product410_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product410_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product410_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product410_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product410_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product410_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product510_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product510_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product510_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product510_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product510_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product510_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product510_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product610_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product610_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product710_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product710_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product710_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product710_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product710_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product710_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product710_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product810_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product810_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product910_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product910_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product910_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product910_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product910_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product910_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product910_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No144_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No145_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No146_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No147_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No148_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No149_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No150_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No151_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No152_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No153_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No154_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No155_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No156_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No157_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No158_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No159_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No160_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No161_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No162_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No163_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No164_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No165_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No166_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No167_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No168_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No169_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No170_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No171_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No172_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No173_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No174_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No175_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No176_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No177_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No178_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No179_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No180_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No181_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No182_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No183_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No184_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No185_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No186_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No187_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No188_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No189_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No190_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No191_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No192_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No193_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No194_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No195_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No196_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No197_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No198_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No199_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No200_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No201_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No202_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No203_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No204_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No205_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No206_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No207_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No208_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No209_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No210_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No211_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No212_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No213_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No214_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No215_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No216_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add30_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add30_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add110_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add110_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add110_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add110_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add110_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add101_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add101_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add101_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add101_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add111_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add111_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add111_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add141_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add141_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add141_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add141_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add141_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add141_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add141_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add141_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add141_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add141_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add141_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add141_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add151_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add151_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No254_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add151_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No255_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add21_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add21_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No256_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add21_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No257_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add23_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add23_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No258_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add23_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No259_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product312_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product312_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No260_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product312_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No261_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product312_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product312_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No262_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product312_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No263_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product312_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product312_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No264_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product312_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No265_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product312_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product312_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No266_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product312_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No267_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product312_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product312_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No268_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product312_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No269_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product312_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product312_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No270_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product312_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No271_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product54_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product54_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No272_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product54_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No273_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product54_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product54_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No274_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product54_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No275_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product62_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product62_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No276_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product62_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No277_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No278_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No279_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No280_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No281_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No282_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No283_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No284_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No285_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_4_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_4_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No286_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_4_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No287_out : std_logic_vector(33 downto 0) := (others => '0');
signal Subtract12_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No288_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Subtract12_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No289_out : std_logic_vector(33 downto 0) := (others => '0');
signal Add10_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add10_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No290_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add10_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No291_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Divide_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Divide_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No292_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Divide_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No293_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product213_5_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_5_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No294_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product213_5_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No295_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No332_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No333_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No334_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No335_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No336_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No337_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No338_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No339_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No340_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No341_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No342_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No343_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No344_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No345_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No346_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No347_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No348_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No349_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay58No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No22_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No39_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay62No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay67No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay24No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay24No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No20_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay59No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay89No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay89No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay69No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay69No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay70No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay70No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay70No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay70No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay70No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay70No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay60No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay60No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay60No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay60No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay55No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay55No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay55No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay55No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay69No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay20No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay48No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay48No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No26_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No24_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No25_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No27_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No29_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Add141_5_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Add141_5_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product62_5_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product62_5_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Add10_5_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Add10_5_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Divide_0_impl_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Divide_0_impl_1_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Product213_5_impl_0_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal MUX_Product213_5_impl_1_LUT_out : std_logic_vector(3 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg581_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg618_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg735_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg959_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg970_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg988_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg989_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg992_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg995_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg996_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1019_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1035_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1040_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1041_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1045_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1048_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1053_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1071_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1074_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1083_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out : std_logic_vector(33 downto 0) := (others => '0');
signal Ldiff_UU_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UU_del_1_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UU_del_1_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UU_del_1_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UU_del_1_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UU_del_1_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UV_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UV_del_1_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UV_del_1_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UV_del_1_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UV_del_1_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UV_del_1_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UW_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UW_del_1_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UW_del_1_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UW_del_1_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UW_del_1_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_UW_del_1_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VU_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VU_del_1_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VU_del_1_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VU_del_1_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VU_del_1_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VU_del_1_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VV_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VV_del_1_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VV_del_1_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VV_del_1_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VV_del_1_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VV_del_1_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VW_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VW_del_1_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VW_del_1_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VW_del_1_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VW_del_1_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_VW_del_1_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WU_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WU_del_1_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WU_del_1_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WU_del_1_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WU_del_1_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WU_del_1_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WV_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WV_del_1_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WV_del_1_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WV_del_1_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WV_del_1_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WV_del_1_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WW_del_1_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WW_del_1_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WW_del_1_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WW_del_1_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WW_del_1_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Ldiff_WW_del_1_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_U_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_U_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_U_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_U_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_U_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_U_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_V_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_V_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_V_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_V_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_V_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_V_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_W_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_W_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_W_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_W_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_W_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal R_W_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Delay1No_out_to_Product108_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out_to_Product108_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1300_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg451_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg779_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg361_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1300_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg927_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No12_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1311_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No6_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out_to_Product108_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out_to_Product108_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No344_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg775_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg542_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg787_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg368_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg981_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No13_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg996_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1311_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out_to_Product108_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out_to_Product108_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No339_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg840_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg553_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg847_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg421_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg992_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1297_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg995_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No14_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out_to_Product108_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out_to_Product108_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg844_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg431_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg849_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1297_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1006_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No15_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out_to_Product108_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out_to_Product108_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No3_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1101_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg860_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1292_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1311_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1297_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1014_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out_to_Product108_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out_to_Product108_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1177_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1193_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1177_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No336_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1199_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg972_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1121_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1116_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1285_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out_to_Product110_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out_to_Product110_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1315_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1302_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg682_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1315_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1302_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg982_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1294_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out_to_Product110_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out_to_Product110_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg364_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1300_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1302_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg638_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg789_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg503_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No7_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1300_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1302_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No1_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg996_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1294_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out_to_Product110_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out_to_Product110_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg372_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No345_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg376_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg785_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1302_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg644_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg647_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1311_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No8_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1302_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No2_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1007_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out_to_Product110_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out_to_Product110_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg856_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg429_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No334_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg384_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg794_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1302_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1302_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No3_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No20_out_to_Product110_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No21_out_to_Product110_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg712_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1197_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No335_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg393_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg855_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No16_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1029_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1285_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No22_out_to_Product110_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No23_out_to_Product110_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1315_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1181_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No342_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1315_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No17_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1294_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1311_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1314_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1289_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No24_out_to_Product109_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No25_out_to_Product109_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg405_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg455_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg727_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1307_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1139_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1310_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No26_out_to_Product109_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No27_out_to_Product109_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg417_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg786_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No1_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1289_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1310_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No28_out_to_Product109_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No29_out_to_Product109_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg797_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No8_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg836_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg784_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1294_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No2_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1314_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1289_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1129_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No30_out_to_Product109_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No31_out_to_Product109_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg803_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg805_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No340_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg895_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg653_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1098_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1294_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1311_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1314_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1289_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg967_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No32_out_to_Product109_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No33_out_to_Product109_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1302_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg663_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg570_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg441_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No341_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1169_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg662_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1302_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No4_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1314_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1289_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No34_out_to_Product109_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No35_out_to_Product109_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg625_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1302_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1192_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No348_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1300_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1046_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1302_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1300_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No36_out_to_Product111_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No37_out_to_Product111_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1313_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg679_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay62No_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg537_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1312_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1313_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1312_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1089_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No38_out_to_Product111_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No39_out_to_Product111_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1313_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1315_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg737_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg462_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg546_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1313_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1315_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No40_out_to_Product111_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No41_out_to_Product111_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg846_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1300_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1315_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg750_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg467_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg555_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1310_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1300_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1315_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No42_out_to_Product111_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No43_out_to_Product111_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1172_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No346_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1300_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1315_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg903_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1310_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1300_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1315_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No44_out_to_Product111_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No45_out_to_Product111_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg813_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg853_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No347_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1300_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1315_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg973_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1300_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1315_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No46_out_to_Product111_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No47_out_to_Product111_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1187_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg527_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg872_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1251_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1311_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No11_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1107_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No48_out_to_Product210_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No49_out_to_Product210_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg495_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1293_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg539_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg940_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1293_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1144_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg984_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No50_out_to_Product210_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No51_out_to_Product210_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1312_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg461_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg366_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1293_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1312_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg941_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg951_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1293_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1066_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No52_out_to_Product210_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No53_out_to_Product210_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1312_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg464_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg509_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1293_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1312_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1020_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1293_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No54_out_to_Product210_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No55_out_to_Product210_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg516_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg562_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg560_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No9_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1031_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1100_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No56_out_to_Product210_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No57_out_to_Product210_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg523_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg863_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg434_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg521_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1270_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1311_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No10_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1118_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1077_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No58_out_to_Product210_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No59_out_to_Product210_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg529_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg620_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg619_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg725_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No11_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1307_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1052_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1308_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay97No5_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1251_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1294_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No5_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No60_out_to_Product310_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No61_out_to_Product310_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg536_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg402_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg497_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg538_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1087_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No62_out_to_Product310_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No63_out_to_Product310_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No7_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg545_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg549_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg457_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg547_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg596_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg997_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1307_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg938_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No64_out_to_Product310_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No65_out_to_Product310_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg556_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg506_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg650_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg698_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1025_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg952_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1307_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg948_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No66_out_to_Product310_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No67_out_to_Product310_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1293_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No9_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg564_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg652_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg659_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1293_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1039_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No3_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1307_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1133_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No68_out_to_Product310_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No69_out_to_Product310_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg666_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg519_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg614_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg816_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay87No10_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg572_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1294_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay102No4_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1307_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No70_out_to_Product310_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No71_out_to_Product310_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg877_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1313_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No5_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1267_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1268_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1269_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1310_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1053_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1313_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No72_out_to_Product410_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No73_out_to_Product410_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No18_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg493_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg588_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1141_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No24_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No74_out_to_Product410_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No75_out_to_Product410_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No19_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg736_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg499_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg992_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1063_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No25_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No76_out_to_Product410_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No77_out_to_Product410_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg651_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1313_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No20_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg793_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg792_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1008_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1313_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1022_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No78_out_to_Product410_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No79_out_to_Product410_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg707_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1313_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg861_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg902_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1313_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay9No39_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No80_out_to_Product410_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No81_out_to_Product410_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1293_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1178_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1313_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1075_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1293_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1310_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1271_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1299_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1273_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1313_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1265_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1119_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No82_out_to_Product410_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No83_out_to_Product410_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg875_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg626_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg623_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1312_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg577_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1109_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1312_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1252_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No84_out_to_Product510_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No85_out_to_Product510_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg776_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg830_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No6_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg932_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1316_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1304_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg990_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No86_out_to_Product510_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No87_out_to_Product510_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg640_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg783_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg838_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg411_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No7_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No1_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1068_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1316_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1304_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No88_out_to_Product510_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No89_out_to_Product510_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg504_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg696_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg552_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg694_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1161_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg646_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg381_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg955_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1003_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No2_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg963_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1316_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1304_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No90_out_to_Product510_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No91_out_to_Product510_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg801_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1312_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg704_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No27_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1312_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1135_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No3_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1041_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1316_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No92_out_to_Product510_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No93_out_to_Product510_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg870_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg909_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg810_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg717_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1312_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg661_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1312_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1078_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay94No4_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1079_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No94_out_to_Product510_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No95_out_to_Product510_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg718_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg826_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg621_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg490_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1293_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg673_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1056_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1293_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1112_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No96_out_to_Product610_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No97_out_to_Product610_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg629_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg677_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg630_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg731_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg452_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg535_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg728_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg929_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1298_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1145_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No98_out_to_Product610_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No99_out_to_Product610_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No1_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No1_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg637_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg743_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg501_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg544_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1001_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg985_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1298_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No100_out_to_Product610_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No101_out_to_Product610_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg508_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No2_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg697_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg597_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg746_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg693_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg753_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg998_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1298_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No102_out_to_Product610_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No103_out_to_Product610_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg390_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg514_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg660_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg706_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg852_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg758_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg807_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1304_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1099_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg961_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1298_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No104_out_to_Product610_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No105_out_to_Product610_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg812_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No10_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg715_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg709_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1316_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1123_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg974_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1036_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No106_out_to_Product610_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No107_out_to_Product610_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg873_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg914_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg674_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1015_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1316_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1050_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No108_out_to_Product710_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No109_out_to_Product710_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1085_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1090_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg777_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg729_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg986_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg979_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg926_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1146_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1296_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1142_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No110_out_to_Product710_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No111_out_to_Product710_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg739_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg942_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg837_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg740_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1067_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg945_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1069_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1296_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1064_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No112_out_to_Product710_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No113_out_to_Product710_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg604_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg900_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No2_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg947_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg954_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg896_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg845_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1010_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg958_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1027_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1296_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1023_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No114_out_to_Product710_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No115_out_to_Product710_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg607_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg657_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1132_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1136_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg389_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1030_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1043_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1296_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No116_out_to_Product710_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No117_out_to_Product710_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg865_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg869_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg612_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1195_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1074_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1298_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1304_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1306_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1287_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No118_out_to_Product710_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No119_out_to_Product710_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg770_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No5_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1317_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No29_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1254_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No11_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No120_out_to_Product810_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No121_out_to_Product810_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg781_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg832_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg831_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1088_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1301_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1291_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1143_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1138_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1285_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No122_out_to_Product810_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No123_out_to_Product810_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg999_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg839_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg891_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg939_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1157_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1019_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1291_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1065_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No124_out_to_Product810_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No125_out_to_Product810_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg796_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg897_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg748_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg791_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg899_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg898_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg949_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1026_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No8_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1291_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No126_out_to_Product810_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No127_out_to_Product810_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg854_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg804_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg802_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg800_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg904_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1033_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No9_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1291_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No128_out_to_Product810_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No129_out_to_Product810_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1080_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1194_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg864_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg814_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg908_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1125_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1296_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1081_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay78No10_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1264_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1117_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No130_out_to_Product810_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No131_out_to_Product810_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1190_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1058_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg773_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1186_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg491_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No5_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1301_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg969_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1114_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1304_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1113_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No132_out_to_Product910_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No133_out_to_Product910_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No332_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg833_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg834_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1149_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg730_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg414_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1297_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg925_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1290_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1303_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1294_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1311_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No134_out_to_Product910_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No135_out_to_Product910_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg636_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1154_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg373_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg741_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg842_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1285_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1060_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1290_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1303_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1294_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1311_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No136_out_to_Product910_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No137_out_to_Product910_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1164_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1009_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg645_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg472_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg512_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg752_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1024_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1018_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1290_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1303_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No138_out_to_Product910_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No139_out_to_Product910_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg438_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1134_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg858_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No3_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No3_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg703_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg518_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1034_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1103_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1128_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1290_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No140_out_to_Product910_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No141_out_to_Product910_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg809_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg399_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg520_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay80No4_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay90No4_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1291_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1120_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg976_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1286_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1277_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg966_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No142_out_to_Product910_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No143_out_to_Product910_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1048_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1256_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg921_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg575_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg723_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg878_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1253_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1258_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1250_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1297_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1012_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1298_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Inv_11_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_11_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_11_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_11_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_11_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_11_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_12_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_12_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_12_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_12_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_12_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_12_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_13_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_13_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_13_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_13_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_13_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_13_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_21_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_21_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_21_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_21_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_21_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_21_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_22_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_22_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_22_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_22_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_22_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_22_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_23_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_23_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_23_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_23_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_23_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_23_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_31_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_31_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_31_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_31_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_31_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_31_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_32_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_32_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_32_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_32_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_32_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_32_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_33_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_33_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_33_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_33_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_33_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_33_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_41_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_41_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_41_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_41_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_41_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_41_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_42_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_42_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_42_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_42_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_42_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_42_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_43_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_43_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_43_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_43_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_43_4_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Inv_43_5_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Delay1No216_out_to_Add30_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No217_out_to_Add30_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg633_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg585_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg403_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg886_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg582_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg450_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg498_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No6_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No6_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg930_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg583_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg531_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay70No_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg584_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No218_out_to_Add30_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No219_out_to_Add30_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg369_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg416_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg502_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1155_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg456_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg459_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg639_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No1_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No1_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg422_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg885_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg532_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No1_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg589_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg641_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No220_out_to_Add30_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No221_out_to_Add30_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg738_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg541_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg466_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg470_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg463_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg554_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg648_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No2_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg841_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg548_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1156_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1000_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg599_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No2_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg642_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg425_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1221_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No222_out_to_Add30_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No223_out_to_Add30_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay24No2_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No8_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg551_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg608_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg605_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg561_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg656_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1163_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1227_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg423_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1037_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg654_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No3_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg755_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg598_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No224_out_to_Add30_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No225_out_to_Add30_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg437_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay60No3_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg808_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg485_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No3_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No10_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1182_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay69No10_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg445_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1198_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg571_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg436_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg957_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1234_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1097_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1236_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No226_out_to_Add30_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No227_out_to_Add30_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No16_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg528_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1211_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay60No4_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay89No10_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1180_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1175_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No11_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1262_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg670_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg448_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg669_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay70No5_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1071_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg398_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1244_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No228_out_to_Add110_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No229_out_to_Add110_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg627_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg593_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay55No6_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No12_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg410_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay19No13_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg540_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay69No12_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg494_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg404_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1220_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg987_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg591_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay70No1_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg887_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg592_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg590_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg359_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No230_out_to_Add110_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No231_out_to_Add110_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg415_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg500_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg634_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg600_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg375_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1158_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay55No7_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No13_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1166_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg747_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg594_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg458_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg413_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg418_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay70No2_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No232_out_to_Add110_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No233_out_to_Add110_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg892_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg888_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg469_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg505_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg699_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg385_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg383_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1165_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay55No8_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No14_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg559_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No2_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg745_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg602_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg465_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg511_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay70No3_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg934_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No234_out_to_Add110_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No235_out_to_Add110_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg446_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg763_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg906_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1168_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg616_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg567_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No11_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg672_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg568_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg764_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg613_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg481_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay67No4_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg971_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1244_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay70No4_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No236_out_to_Add101_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No237_out_to_Add101_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg468_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No1_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No8_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg799_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg507_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1162_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg692_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg603_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No8_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1163_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No7_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1222_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1224_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1226_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg754_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1225_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg471_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg749_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No238_out_to_Add101_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No239_out_to_Add101_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg563_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No9_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No3_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg558_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg664_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg768_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg665_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No9_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg756_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay6No3_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg474_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg476_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1238_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1016_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No4_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No240_out_to_Add101_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No241_out_to_Add101_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg526_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg823_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No5_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg487_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg675_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg923_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1210_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg719_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay69No11_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg772_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay96No5_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg720_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg525_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1247_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1045_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg771_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No242_out_to_Add111_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No243_out_to_Add111_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No7_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No7_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg689_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1159_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg686_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg365_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg595_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No7_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg889_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1153_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg890_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay24No1_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg937_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1218_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg744_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1219_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg371_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1223_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1216_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No244_out_to_Add111_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No245_out_to_Add111_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No4_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No4_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay14No4_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg615_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No10_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg766_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg611_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg447_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg579_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg580_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1196_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg714_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg716_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1241_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1176_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg576_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1239_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No246_out_to_Add141_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No247_out_to_Add141_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg496_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1150_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg678_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg631_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg412_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No6_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg406_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg407_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1214_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg732_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1215_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg879_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg632_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg363_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1217_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg453_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No248_out_to_Add141_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No249_out_to_Add141_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1160_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No8_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg477_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No2_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg475_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg478_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg513_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg388_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg757_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg473_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg655_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1173_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg430_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg379_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1229_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1228_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1232_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg761_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg649_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No250_out_to_Add141_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No251_out_to_Add141_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No3_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg440_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1167_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No9_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg606_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg483_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg617_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg569_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg395_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg811_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No15_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg479_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1231_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg658_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg386_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1235_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1170_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1233_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1238_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg817_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg517_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1127_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No252_out_to_Add141_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No253_out_to_Add141_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No11_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No5_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay104No5_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg774_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg819_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1209_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg874_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1260_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg578_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg724_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg825_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1246_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1243_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1207_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No254_out_to_Add151_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No255_out_to_Add151_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No10_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg396_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1174_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg397_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1191_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg449_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg818_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No11_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg722_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg922_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay59No5_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg667_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg442_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1094_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg394_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1241_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1240_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1245_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1054_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1237_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No256_out_to_Add21_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No257_out_to_Add21_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg850_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay89No8_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No26_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg894_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay88No9_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay76No9_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg708_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg482_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg392_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg391_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg484_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No3_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg428_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg944_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1230_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1230_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg433_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No258_out_to_Add23_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No259_out_to_Add23_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg683_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg884_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg883_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1152_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No6_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg829_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg827_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg882_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay60No_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg734_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg586_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg733_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1213_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1148_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1082_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1083_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1151_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1212_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No260_out_to_Product312_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No261_out_to_Product312_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No338_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg880_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg778_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg400_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg681_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg726_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg881_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg828_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1314_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1292_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1137_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg978_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No262_out_to_Product312_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No263_out_to_Product312_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg424_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No333_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg936_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg790_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg408_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg782_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg742_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg835_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg420_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg993_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1301_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1292_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1059_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No264_out_to_Product312_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No265_out_to_Product312_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg851_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1162_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg380_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg946_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg798_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg550_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg893_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg848_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg843_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg427_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1294_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1311_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1285_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1005_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1301_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1292_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No266_out_to_Product312_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No267_out_to_Product312_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg760_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg435_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1171_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg905_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg387_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1131_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg806_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg557_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg901_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg859_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1303_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1294_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1040_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1096_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1301_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No268_out_to_Product312_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No269_out_to_Product312_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg443_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg489_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg815_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1076_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg767_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1070_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg912_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg488_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1073_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg868_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg566_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1290_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1303_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1282_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1124_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1275_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg970_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1301_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No270_out_to_Product312_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No271_out_to_Product312_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1186_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg524_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg916_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg821_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg919_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg822_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1290_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1296_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1309_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1110_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1285_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No272_out_to_Product54_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No273_out_to_Product54_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg907_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg867_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg862_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1179_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg910_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg975_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay20No16_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg610_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1292_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1297_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No274_out_to_Product54_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No275_out_to_Product54_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1189_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg573_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1204_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1203_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1051_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg917_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1262_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1186_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No337_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1276_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1288_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1291_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1280_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1111_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1283_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1105_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1305_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1295_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No276_out_to_Product62_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No277_out_to_Product62_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No343_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1184_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1200_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg920_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay64No5_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1259_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg913_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1249_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1314_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1278_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1311_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1294_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1284_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1303_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No278_out_to_Subtract12_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No279_out_to_Subtract12_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg587_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg454_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg360_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg534_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg680_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg780_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg362_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg533_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg676_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay48No_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg401_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg628_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay73No_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1086_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1084_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1147_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg931_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg928_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1140_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg980_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg924_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No280_out_to_Subtract12_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No281_out_to_Subtract12_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg409_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg635_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg688_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg460_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No1_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg367_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg543_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg687_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg788_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg370_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg685_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg684_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg377_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg994_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg989_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1062_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg935_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No1_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg988_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg983_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg933_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1061_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No282_out_to_Subtract12_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No283_out_to_Subtract12_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg690_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay48No2_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg419_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg643_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg695_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg510_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No2_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg374_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg601_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg751_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg795_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg378_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg691_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1004_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg991_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg959_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg953_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1021_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1092_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No2_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1002_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg962_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg950_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg943_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No284_out_to_Subtract12_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No285_out_to_Subtract12_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg432_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg702_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg700_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg522_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg426_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg701_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg705_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg515_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg565_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg382_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg609_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg759_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg857_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg956_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1130_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1032_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg964_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1093_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1095_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1102_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1038_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg960_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No286_out_to_Subtract12_4_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No287_out_to_Subtract12_4_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg911_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg866_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg486_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg711_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg762_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg492_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg480_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg710_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg713_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg668_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No4_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg439_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg765_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay58No4_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1035_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1028_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No22_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1042_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1013_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1072_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay79No4_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1011_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No288_out_to_Subtract12_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No289_out_to_Subtract12_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay84No5_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg444_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg721_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg876_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1188_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg530_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg671_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1261_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg574_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg820_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg622_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg624_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1106_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1126_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1055_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1122_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1047_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1108_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1044_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1057_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1049_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No290_out_to_Add10_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No291_out_to_Add10_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay5No17_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay60No5_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay55No11_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg871_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg918_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1206_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1202_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1205_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1242_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1257_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No292_out_to_Divide_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No293_out_to_Divide_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1255_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg977_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1017_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1091_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg965_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1115_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg968_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No294_out_to_Product213_5_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No295_out_to_Product213_5_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No349_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg915_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1185_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1201_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg769_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1208_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg824_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1183_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1248_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1104_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1274_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1279_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1281_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1266_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1292_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1272_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1289_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1263_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount131_instance: ModuloCounter_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount131_out);
Ldiff_UU_del_1_0_IEEE <= Ldiff_UU_del_1_0;
   Ldiff_UU_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UU_del_1_0_out,
                 X => Ldiff_UU_del_1_0_IEEE);
Ldiff_UU_del_1_1_IEEE <= Ldiff_UU_del_1_1;
   Ldiff_UU_del_1_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UU_del_1_1_out,
                 X => Ldiff_UU_del_1_1_IEEE);
Ldiff_UU_del_1_2_IEEE <= Ldiff_UU_del_1_2;
   Ldiff_UU_del_1_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UU_del_1_2_out,
                 X => Ldiff_UU_del_1_2_IEEE);
Ldiff_UU_del_1_3_IEEE <= Ldiff_UU_del_1_3;
   Ldiff_UU_del_1_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UU_del_1_3_out,
                 X => Ldiff_UU_del_1_3_IEEE);
Ldiff_UU_del_1_4_IEEE <= Ldiff_UU_del_1_4;
   Ldiff_UU_del_1_4_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UU_del_1_4_out,
                 X => Ldiff_UU_del_1_4_IEEE);
Ldiff_UU_del_1_5_IEEE <= Ldiff_UU_del_1_5;
   Ldiff_UU_del_1_5_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UU_del_1_5_out,
                 X => Ldiff_UU_del_1_5_IEEE);
Ldiff_UV_del_1_0_IEEE <= Ldiff_UV_del_1_0;
   Ldiff_UV_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UV_del_1_0_out,
                 X => Ldiff_UV_del_1_0_IEEE);
Ldiff_UV_del_1_1_IEEE <= Ldiff_UV_del_1_1;
   Ldiff_UV_del_1_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UV_del_1_1_out,
                 X => Ldiff_UV_del_1_1_IEEE);
Ldiff_UV_del_1_2_IEEE <= Ldiff_UV_del_1_2;
   Ldiff_UV_del_1_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UV_del_1_2_out,
                 X => Ldiff_UV_del_1_2_IEEE);
Ldiff_UV_del_1_3_IEEE <= Ldiff_UV_del_1_3;
   Ldiff_UV_del_1_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UV_del_1_3_out,
                 X => Ldiff_UV_del_1_3_IEEE);
Ldiff_UV_del_1_4_IEEE <= Ldiff_UV_del_1_4;
   Ldiff_UV_del_1_4_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UV_del_1_4_out,
                 X => Ldiff_UV_del_1_4_IEEE);
Ldiff_UV_del_1_5_IEEE <= Ldiff_UV_del_1_5;
   Ldiff_UV_del_1_5_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UV_del_1_5_out,
                 X => Ldiff_UV_del_1_5_IEEE);
Ldiff_UW_del_1_0_IEEE <= Ldiff_UW_del_1_0;
   Ldiff_UW_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UW_del_1_0_out,
                 X => Ldiff_UW_del_1_0_IEEE);
Ldiff_UW_del_1_1_IEEE <= Ldiff_UW_del_1_1;
   Ldiff_UW_del_1_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UW_del_1_1_out,
                 X => Ldiff_UW_del_1_1_IEEE);
Ldiff_UW_del_1_2_IEEE <= Ldiff_UW_del_1_2;
   Ldiff_UW_del_1_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UW_del_1_2_out,
                 X => Ldiff_UW_del_1_2_IEEE);
Ldiff_UW_del_1_3_IEEE <= Ldiff_UW_del_1_3;
   Ldiff_UW_del_1_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UW_del_1_3_out,
                 X => Ldiff_UW_del_1_3_IEEE);
Ldiff_UW_del_1_4_IEEE <= Ldiff_UW_del_1_4;
   Ldiff_UW_del_1_4_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UW_del_1_4_out,
                 X => Ldiff_UW_del_1_4_IEEE);
Ldiff_UW_del_1_5_IEEE <= Ldiff_UW_del_1_5;
   Ldiff_UW_del_1_5_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_UW_del_1_5_out,
                 X => Ldiff_UW_del_1_5_IEEE);
Ldiff_VU_del_1_0_IEEE <= Ldiff_VU_del_1_0;
   Ldiff_VU_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VU_del_1_0_out,
                 X => Ldiff_VU_del_1_0_IEEE);
Ldiff_VU_del_1_1_IEEE <= Ldiff_VU_del_1_1;
   Ldiff_VU_del_1_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VU_del_1_1_out,
                 X => Ldiff_VU_del_1_1_IEEE);
Ldiff_VU_del_1_2_IEEE <= Ldiff_VU_del_1_2;
   Ldiff_VU_del_1_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VU_del_1_2_out,
                 X => Ldiff_VU_del_1_2_IEEE);
Ldiff_VU_del_1_3_IEEE <= Ldiff_VU_del_1_3;
   Ldiff_VU_del_1_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VU_del_1_3_out,
                 X => Ldiff_VU_del_1_3_IEEE);
Ldiff_VU_del_1_4_IEEE <= Ldiff_VU_del_1_4;
   Ldiff_VU_del_1_4_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VU_del_1_4_out,
                 X => Ldiff_VU_del_1_4_IEEE);
Ldiff_VU_del_1_5_IEEE <= Ldiff_VU_del_1_5;
   Ldiff_VU_del_1_5_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VU_del_1_5_out,
                 X => Ldiff_VU_del_1_5_IEEE);
Ldiff_VV_del_1_0_IEEE <= Ldiff_VV_del_1_0;
   Ldiff_VV_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VV_del_1_0_out,
                 X => Ldiff_VV_del_1_0_IEEE);
Ldiff_VV_del_1_1_IEEE <= Ldiff_VV_del_1_1;
   Ldiff_VV_del_1_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VV_del_1_1_out,
                 X => Ldiff_VV_del_1_1_IEEE);
Ldiff_VV_del_1_2_IEEE <= Ldiff_VV_del_1_2;
   Ldiff_VV_del_1_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VV_del_1_2_out,
                 X => Ldiff_VV_del_1_2_IEEE);
Ldiff_VV_del_1_3_IEEE <= Ldiff_VV_del_1_3;
   Ldiff_VV_del_1_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VV_del_1_3_out,
                 X => Ldiff_VV_del_1_3_IEEE);
Ldiff_VV_del_1_4_IEEE <= Ldiff_VV_del_1_4;
   Ldiff_VV_del_1_4_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VV_del_1_4_out,
                 X => Ldiff_VV_del_1_4_IEEE);
Ldiff_VV_del_1_5_IEEE <= Ldiff_VV_del_1_5;
   Ldiff_VV_del_1_5_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VV_del_1_5_out,
                 X => Ldiff_VV_del_1_5_IEEE);
Ldiff_VW_del_1_0_IEEE <= Ldiff_VW_del_1_0;
   Ldiff_VW_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VW_del_1_0_out,
                 X => Ldiff_VW_del_1_0_IEEE);
Ldiff_VW_del_1_1_IEEE <= Ldiff_VW_del_1_1;
   Ldiff_VW_del_1_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VW_del_1_1_out,
                 X => Ldiff_VW_del_1_1_IEEE);
Ldiff_VW_del_1_2_IEEE <= Ldiff_VW_del_1_2;
   Ldiff_VW_del_1_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VW_del_1_2_out,
                 X => Ldiff_VW_del_1_2_IEEE);
Ldiff_VW_del_1_3_IEEE <= Ldiff_VW_del_1_3;
   Ldiff_VW_del_1_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VW_del_1_3_out,
                 X => Ldiff_VW_del_1_3_IEEE);
Ldiff_VW_del_1_4_IEEE <= Ldiff_VW_del_1_4;
   Ldiff_VW_del_1_4_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VW_del_1_4_out,
                 X => Ldiff_VW_del_1_4_IEEE);
Ldiff_VW_del_1_5_IEEE <= Ldiff_VW_del_1_5;
   Ldiff_VW_del_1_5_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_VW_del_1_5_out,
                 X => Ldiff_VW_del_1_5_IEEE);
Ldiff_WU_del_1_0_IEEE <= Ldiff_WU_del_1_0;
   Ldiff_WU_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WU_del_1_0_out,
                 X => Ldiff_WU_del_1_0_IEEE);
Ldiff_WU_del_1_1_IEEE <= Ldiff_WU_del_1_1;
   Ldiff_WU_del_1_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WU_del_1_1_out,
                 X => Ldiff_WU_del_1_1_IEEE);
Ldiff_WU_del_1_2_IEEE <= Ldiff_WU_del_1_2;
   Ldiff_WU_del_1_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WU_del_1_2_out,
                 X => Ldiff_WU_del_1_2_IEEE);
Ldiff_WU_del_1_3_IEEE <= Ldiff_WU_del_1_3;
   Ldiff_WU_del_1_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WU_del_1_3_out,
                 X => Ldiff_WU_del_1_3_IEEE);
Ldiff_WU_del_1_4_IEEE <= Ldiff_WU_del_1_4;
   Ldiff_WU_del_1_4_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WU_del_1_4_out,
                 X => Ldiff_WU_del_1_4_IEEE);
Ldiff_WU_del_1_5_IEEE <= Ldiff_WU_del_1_5;
   Ldiff_WU_del_1_5_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WU_del_1_5_out,
                 X => Ldiff_WU_del_1_5_IEEE);
Ldiff_WV_del_1_0_IEEE <= Ldiff_WV_del_1_0;
   Ldiff_WV_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WV_del_1_0_out,
                 X => Ldiff_WV_del_1_0_IEEE);
Ldiff_WV_del_1_1_IEEE <= Ldiff_WV_del_1_1;
   Ldiff_WV_del_1_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WV_del_1_1_out,
                 X => Ldiff_WV_del_1_1_IEEE);
Ldiff_WV_del_1_2_IEEE <= Ldiff_WV_del_1_2;
   Ldiff_WV_del_1_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WV_del_1_2_out,
                 X => Ldiff_WV_del_1_2_IEEE);
Ldiff_WV_del_1_3_IEEE <= Ldiff_WV_del_1_3;
   Ldiff_WV_del_1_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WV_del_1_3_out,
                 X => Ldiff_WV_del_1_3_IEEE);
Ldiff_WV_del_1_4_IEEE <= Ldiff_WV_del_1_4;
   Ldiff_WV_del_1_4_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WV_del_1_4_out,
                 X => Ldiff_WV_del_1_4_IEEE);
Ldiff_WV_del_1_5_IEEE <= Ldiff_WV_del_1_5;
   Ldiff_WV_del_1_5_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WV_del_1_5_out,
                 X => Ldiff_WV_del_1_5_IEEE);
Ldiff_WW_del_1_0_IEEE <= Ldiff_WW_del_1_0;
   Ldiff_WW_del_1_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WW_del_1_0_out,
                 X => Ldiff_WW_del_1_0_IEEE);
Ldiff_WW_del_1_1_IEEE <= Ldiff_WW_del_1_1;
   Ldiff_WW_del_1_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WW_del_1_1_out,
                 X => Ldiff_WW_del_1_1_IEEE);
Ldiff_WW_del_1_2_IEEE <= Ldiff_WW_del_1_2;
   Ldiff_WW_del_1_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WW_del_1_2_out,
                 X => Ldiff_WW_del_1_2_IEEE);
Ldiff_WW_del_1_3_IEEE <= Ldiff_WW_del_1_3;
   Ldiff_WW_del_1_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WW_del_1_3_out,
                 X => Ldiff_WW_del_1_3_IEEE);
Ldiff_WW_del_1_4_IEEE <= Ldiff_WW_del_1_4;
   Ldiff_WW_del_1_4_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WW_del_1_4_out,
                 X => Ldiff_WW_del_1_4_IEEE);
Ldiff_WW_del_1_5_IEEE <= Ldiff_WW_del_1_5;
   Ldiff_WW_del_1_5_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Ldiff_WW_del_1_5_out,
                 X => Ldiff_WW_del_1_5_IEEE);
R_U_0_IEEE <= R_U_0;
   R_U_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_U_0_out,
                 X => R_U_0_IEEE);
R_U_1_IEEE <= R_U_1;
   R_U_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_U_1_out,
                 X => R_U_1_IEEE);
R_U_2_IEEE <= R_U_2;
   R_U_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_U_2_out,
                 X => R_U_2_IEEE);
R_U_3_IEEE <= R_U_3;
   R_U_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_U_3_out,
                 X => R_U_3_IEEE);
R_U_4_IEEE <= R_U_4;
   R_U_4_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_U_4_out,
                 X => R_U_4_IEEE);
R_U_5_IEEE <= R_U_5;
   R_U_5_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_U_5_out,
                 X => R_U_5_IEEE);
R_V_0_IEEE <= R_V_0;
   R_V_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_V_0_out,
                 X => R_V_0_IEEE);
R_V_1_IEEE <= R_V_1;
   R_V_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_V_1_out,
                 X => R_V_1_IEEE);
R_V_2_IEEE <= R_V_2;
   R_V_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_V_2_out,
                 X => R_V_2_IEEE);
R_V_3_IEEE <= R_V_3;
   R_V_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_V_3_out,
                 X => R_V_3_IEEE);
R_V_4_IEEE <= R_V_4;
   R_V_4_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_V_4_out,
                 X => R_V_4_IEEE);
R_V_5_IEEE <= R_V_5;
   R_V_5_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_V_5_out,
                 X => R_V_5_IEEE);
R_W_0_IEEE <= R_W_0;
   R_W_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_W_0_out,
                 X => R_W_0_IEEE);
R_W_1_IEEE <= R_W_1;
   R_W_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_W_1_out,
                 X => R_W_1_IEEE);
R_W_2_IEEE <= R_W_2;
   R_W_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_W_2_out,
                 X => R_W_2_IEEE);
R_W_3_IEEE <= R_W_3;
   R_W_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_W_3_out,
                 X => R_W_3_IEEE);
R_W_4_IEEE <= R_W_4;
   R_W_4_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_W_4_out,
                 X => R_W_4_IEEE);
R_W_5_IEEE <= R_W_5;
   R_W_5_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_W_5_out,
                 X => R_W_5_IEEE);

Delay1No_out_to_Product108_0_impl_parent_implementedSystem_port_0_cast <= Delay1No_out;
Delay1No1_out_to_Product108_0_impl_parent_implementedSystem_port_1_cast <= Delay1No1_out;
   Product108_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_0_impl_out,
                 X => Delay1No_out_to_Product108_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No1_out_to_Product108_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1306_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1306_out;
SharedReg1300_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1300_out;
SharedReg1_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1_out;
SharedReg451_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg451_out;
SharedReg1256_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1256_out;
SharedReg496_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg496_out;
SharedReg1317_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1317_out;
SharedReg779_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg779_out;
SharedReg361_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg361_out;
SharedReg1270_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1270_out;
SharedReg776_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg776_out;
SharedReg355_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg355_out;
SharedReg1273_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1273_out;
   MUX_Product108_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1306_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1300_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg776_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg355_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1273_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg451_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1256_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg496_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1317_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg779_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg361_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1270_out_to_MUX_Product108_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_0_impl_0_out);

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_0_impl_0_out,
                 Y => Delay1No_out);

SharedReg1306_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1306_out;
SharedReg1300_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1300_out;
SharedReg175_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg175_out;
SharedReg183_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg183_out;
SharedReg927_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg927_out;
Delay87No12_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_6_cast <= Delay87No12_out;
SharedReg1317_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1317_out;
SharedReg1280_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1280_out;
SharedReg982_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg982_out;
SharedReg1270_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1270_out;
SharedReg1311_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1311_out;
Delay102No6_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_12_cast <= Delay102No6_out;
SharedReg1273_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1273_out;
   MUX_Product108_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1306_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1300_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1311_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay102No6_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1273_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg175_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg183_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg927_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay87No12_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1317_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1280_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg982_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1270_out_to_MUX_Product108_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_0_impl_1_out);

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_0_impl_1_out,
                 Y => Delay1No1_out);

Delay1No2_out_to_Product108_1_impl_parent_implementedSystem_port_0_cast <= Delay1No2_out;
Delay1No3_out_to_Product108_1_impl_parent_implementedSystem_port_1_cast <= Delay1No3_out;
   Product108_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_1_impl_out,
                 X => Delay1No2_out_to_Product108_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No3_out_to_Product108_1_impl_parent_implementedSystem_port_1_cast);

SharedReg880_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg880_out;
Delay1No344_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_2_cast <= Delay1No344_out;
SharedReg1306_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1306_out;
SharedReg828_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg828_out;
SharedReg450_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg450_out;
SharedReg775_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg775_out;
SharedReg1256_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1256_out;
SharedReg542_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg542_out;
SharedReg1317_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1317_out;
SharedReg787_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg787_out;
SharedReg368_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg368_out;
SharedReg1270_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1270_out;
SharedReg783_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg783_out;
   MUX_Product108_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg880_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No344_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg368_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1270_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg783_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1306_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg828_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg450_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg775_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1256_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg542_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1317_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg787_out_to_MUX_Product108_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_1_impl_0_out);

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_1_impl_0_out,
                 Y => Delay1No2_out);

SharedReg1274_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1263_out;
SharedReg1306_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1306_out;
SharedReg1288_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1288_out;
SharedReg131_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg131_out;
SharedReg1278_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1278_out;
SharedReg981_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg981_out;
Delay87No13_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_8_cast <= Delay87No13_out;
SharedReg1317_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1317_out;
SharedReg1280_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1280_out;
SharedReg996_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg996_out;
SharedReg1270_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1270_out;
SharedReg1311_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1311_out;
   MUX_Product108_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1274_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1263_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg996_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1270_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1311_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1306_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1288_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg131_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1278_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg981_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay87No13_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1317_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1280_out_to_MUX_Product108_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_1_impl_1_out);

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_1_impl_1_out,
                 Y => Delay1No3_out);

Delay1No4_out_to_Product108_2_impl_parent_implementedSystem_port_0_cast <= Delay1No4_out;
Delay1No5_out_to_Product108_2_impl_parent_implementedSystem_port_1_cast <= Delay1No5_out;
   Product108_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_2_impl_out,
                 X => Delay1No4_out_to_Product108_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No5_out_to_Product108_2_impl_parent_implementedSystem_port_1_cast);

SharedReg836_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg836_out;
SharedReg15_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg15_out;
SharedReg888_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg888_out;
Delay1No339_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_4_cast <= Delay1No339_out;
SharedReg310_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg310_out;
SharedReg840_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg840_out;
SharedReg456_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg456_out;
SharedReg835_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg835_out;
SharedReg1256_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1256_out;
SharedReg553_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg553_out;
SharedReg1317_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1317_out;
SharedReg847_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg847_out;
SharedReg421_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg421_out;
   MUX_Product108_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg836_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg15_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1317_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg847_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg421_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg888_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay1No339_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg310_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg840_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg456_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg835_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1256_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg553_out_to_MUX_Product108_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_2_impl_0_out);

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_2_impl_0_out,
                 Y => Delay1No4_out);

SharedReg1272_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1272_out;
SharedReg992_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg992_out;
SharedReg1274_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1263_out;
SharedReg135_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg135_out;
SharedReg1297_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1297_out;
SharedReg139_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg139_out;
SharedReg1278_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1278_out;
SharedReg995_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg995_out;
Delay87No14_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_10_cast <= Delay87No14_out;
SharedReg1317_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1317_out;
SharedReg1280_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1280_out;
SharedReg1007_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1007_out;
   MUX_Product108_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1272_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg992_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1317_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1280_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1007_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1274_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1263_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg135_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1297_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg139_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1278_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg995_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay87No14_out_to_MUX_Product108_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_2_impl_1_out);

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_2_impl_1_out,
                 Y => Delay1No5_out);

Delay1No6_out_to_Product108_3_impl_parent_implementedSystem_port_0_cast <= Delay1No6_out;
Delay1No7_out_to_Product108_3_impl_parent_implementedSystem_port_1_cast <= Delay1No7_out;
   Product108_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_3_impl_out,
                 X => Delay1No6_out_to_Product108_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No7_out_to_Product108_3_impl_parent_implementedSystem_port_1_cast);

SharedReg261_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg261_out;
SharedReg1002_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1002_out;
SharedReg844_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg844_out;
SharedReg431_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg431_out;
SharedReg30_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg30_out;
SharedReg22_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg22_out;
SharedReg319_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg319_out;
SharedReg849_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg849_out;
SharedReg597_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg597_out;
SharedReg1160_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1160_out;
SharedReg1256_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1256_out;
SharedReg703_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg703_out;
SharedReg1317_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1317_out;
   MUX_Product108_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg261_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1002_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1256_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg703_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1317_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg844_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg431_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg30_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg22_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg319_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg849_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg597_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1160_out_to_MUX_Product108_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_3_impl_0_out);

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_3_impl_0_out,
                 Y => Delay1No6_out);

SharedReg199_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg199_out;
SharedReg1017_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1017_out;
SharedReg1272_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1272_out;
SharedReg1305_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1305_out;
SharedReg265_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg265_out;
SharedReg142_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg142_out;
SharedReg143_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg143_out;
SharedReg1297_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1297_out;
SharedReg147_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg147_out;
SharedReg1278_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1278_out;
SharedReg1006_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1006_out;
Delay87No15_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_12_cast <= Delay87No15_out;
SharedReg1317_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1317_out;
   MUX_Product108_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg199_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1017_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1006_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay87No15_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1317_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1272_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1305_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg265_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg142_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg143_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1297_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg147_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1278_out_to_MUX_Product108_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_3_impl_1_out);

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_3_impl_1_out,
                 Y => Delay1No7_out);

Delay1No8_out_to_Product108_4_impl_parent_implementedSystem_port_0_cast <= Delay1No8_out;
Delay1No9_out_to_Product108_4_impl_parent_implementedSystem_port_1_cast <= Delay1No9_out;
   Product108_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_4_impl_out,
                 X => Delay1No8_out_to_Product108_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No9_out_to_Product108_4_impl_parent_implementedSystem_port_1_cast);

SharedReg852_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg852_out;
SharedReg435_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg435_out;
SharedReg271_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg271_out;
Delay64No3_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_4_cast <= Delay64No3_out;
SharedReg903_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg903_out;
SharedReg1101_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1101_out;
SharedReg41_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg41_out;
SharedReg33_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg33_out;
SharedReg328_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg328_out;
SharedReg860_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg860_out;
SharedReg605_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg605_out;
SharedReg1167_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1167_out;
SharedReg1256_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1256_out;
   MUX_Product108_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg852_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg435_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg605_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1167_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1256_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg271_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay64No3_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg903_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1101_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg41_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg33_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg328_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg860_out_to_MUX_Product108_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_4_impl_0_out);

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_4_impl_0_out,
                 Y => Delay1No8_out);

SharedReg1292_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1292_out;
SharedReg1281_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1281_out;
SharedReg210_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg210_out;
SharedReg1311_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1311_out;
SharedReg1284_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1284_out;
SharedReg157_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg157_out;
SharedReg275_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg275_out;
SharedReg150_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg150_out;
SharedReg151_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg151_out;
SharedReg1297_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1297_out;
SharedReg155_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg155_out;
SharedReg1278_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1278_out;
SharedReg1014_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1014_out;
   MUX_Product108_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1292_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1281_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg155_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1278_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1014_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg210_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1311_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1284_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg157_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg275_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg150_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg151_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1297_out_to_MUX_Product108_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_4_impl_1_out);

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_4_impl_1_out,
                 Y => Delay1No9_out);

Delay1No10_out_to_Product108_5_impl_parent_implementedSystem_port_0_cast <= Delay1No10_out;
Delay1No11_out_to_Product108_5_impl_parent_implementedSystem_port_1_cast <= Delay1No11_out;
   Product108_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product108_5_impl_out,
                 X => Delay1No10_out_to_Product108_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No11_out_to_Product108_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1174_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1174_out;
SharedReg619_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg619_out;
SharedReg1256_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1256_out;
SharedReg395_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg395_out;
SharedReg283_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg283_out;
SharedReg1177_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1177_out;
SharedReg110_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg110_out;
SharedReg1193_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1193_out;
SharedReg1177_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1177_out;
Delay1No336_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_10_cast <= Delay1No336_out;
SharedReg1199_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1199_out;
SharedReg910_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg910_out;
SharedReg809_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg809_out;
   MUX_Product108_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1174_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg619_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1199_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg910_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg809_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1256_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg395_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg283_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1177_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg110_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1193_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1177_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay1No336_out_to_MUX_Product108_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_5_impl_0_out);

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_5_impl_0_out,
                 Y => Delay1No10_out);

SharedReg1278_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1278_out;
SharedReg238_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg238_out;
SharedReg972_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg972_out;
SharedReg1281_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1281_out;
SharedReg1121_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1121_out;
SharedReg1283_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1283_out;
SharedReg1116_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1116_out;
SharedReg1285_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1285_out;
SharedReg1295_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1295_out;
SharedReg1263_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1263_out;
SharedReg1276_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1276_out;
SharedReg1288_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1288_out;
SharedReg54_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg54_out;
   MUX_Product108_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1278_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg238_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1276_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1288_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg54_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg972_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1281_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1121_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1283_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1116_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1285_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1295_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1263_out_to_MUX_Product108_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product108_5_impl_1_out);

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product108_5_impl_1_out,
                 Y => Delay1No11_out);

Delay1No12_out_to_Product110_0_impl_parent_implementedSystem_port_0_cast <= Delay1No12_out;
Delay1No13_out_to_Product110_0_impl_parent_implementedSystem_port_1_cast <= Delay1No13_out;
   Product110_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_0_impl_out,
                 X => Delay1No12_out_to_Product110_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No13_out_to_Product110_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1274_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1274_out;
SharedReg452_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg452_out;
SharedReg67_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg67_out;
SharedReg1315_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1315_out;
SharedReg1256_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1256_out;
SharedReg1302_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1302_out;
SharedReg495_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg495_out;
SharedReg494_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg494_out;
SharedReg587_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg587_out;
SharedReg682_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg682_out;
SharedReg358_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg358_out;
SharedReg362_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg362_out;
SharedReg1305_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1305_out;
   MUX_Product110_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1274_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg452_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg358_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg362_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1305_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg67_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1315_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1256_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1302_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg495_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg494_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg587_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg682_out_to_MUX_Product110_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_0_impl_0_out);

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_0_impl_0_out,
                 Y => Delay1No12_out);

SharedReg1274_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1274_out;
SharedReg1140_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1140_out;
SharedReg127_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg127_out;
SharedReg1315_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1315_out;
SharedReg1137_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1137_out;
SharedReg1302_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1302_out;
Delay97No_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_7_cast <= Delay97No_out;
SharedReg302_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg302_out;
SharedReg982_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg982_out;
SharedReg1294_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1294_out;
SharedReg1271_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1271_out;
Delay102No_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_12_cast <= Delay102No_out;
SharedReg1305_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1305_out;
   MUX_Product110_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1274_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1140_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1271_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay102No_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1305_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg127_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1315_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1137_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1302_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay97No_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg302_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg982_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1294_out_to_MUX_Product110_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_0_impl_1_out);

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_0_impl_1_out,
                 Y => Delay1No13_out);

Delay1No14_out_to_Product110_1_impl_parent_implementedSystem_port_0_cast <= Delay1No14_out;
Delay1No15_out_to_Product110_1_impl_parent_implementedSystem_port_1_cast <= Delay1No15_out;
   Product110_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_1_impl_out,
                 X => Delay1No14_out_to_Product110_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No15_out_to_Product110_1_impl_parent_implementedSystem_port_1_cast);

SharedReg364_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg364_out;
SharedReg1273_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1273_out;
SharedReg1274_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1274_out;
SharedReg1300_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1300_out;
SharedReg627_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg627_out;
SharedReg827_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg827_out;
SharedReg1256_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1256_out;
SharedReg1302_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1302_out;
SharedReg501_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg501_out;
SharedReg635_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg635_out;
SharedReg638_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg638_out;
SharedReg789_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg789_out;
SharedReg503_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg503_out;
   MUX_Product110_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg364_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1273_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg638_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg789_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg503_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1274_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1300_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg627_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg827_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1256_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1302_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg501_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg635_out_to_MUX_Product110_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_1_impl_0_out);

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_1_impl_0_out,
                 Y => Delay1No14_out);

Delay102No7_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_1_cast <= Delay102No7_out;
SharedReg1273_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1273_out;
SharedReg1274_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1274_out;
SharedReg1300_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1300_out;
SharedReg10_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg10_out;
SharedReg1266_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1266_out;
SharedReg1059_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1059_out;
SharedReg1302_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1302_out;
Delay97No1_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_9_cast <= Delay97No1_out;
SharedReg311_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg311_out;
SharedReg996_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg996_out;
SharedReg1294_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1294_out;
SharedReg1271_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1271_out;
   MUX_Product110_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay102No7_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1273_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg996_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1294_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1271_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1274_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1300_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg10_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1266_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1059_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1302_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay97No1_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg311_out_to_MUX_Product110_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_1_impl_1_out);

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_1_impl_1_out,
                 Y => Delay1No15_out);

Delay1No16_out_to_Product110_2_impl_parent_implementedSystem_port_0_cast <= Delay1No16_out;
Delay1No17_out_to_Product110_2_impl_parent_implementedSystem_port_1_cast <= Delay1No17_out;
   Product110_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_2_impl_out,
                 X => Delay1No16_out_to_Product110_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No17_out_to_Product110_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1270_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1270_out;
SharedReg792_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg792_out;
SharedReg372_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg372_out;
Delay1No345_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_4_cast <= Delay1No345_out;
SharedReg376_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg376_out;
SharedReg785_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg785_out;
SharedReg634_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg634_out;
SharedReg887_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg887_out;
SharedReg1256_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1256_out;
SharedReg1302_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1302_out;
SharedReg644_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg644_out;
SharedReg643_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg643_out;
SharedReg647_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg647_out;
   MUX_Product110_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1270_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg792_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg644_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg643_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg647_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg372_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay1No345_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg376_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg785_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg634_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg887_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1256_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1302_out_to_MUX_Product110_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_2_impl_0_out);

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_2_impl_0_out,
                 Y => Delay1No16_out);

SharedReg1270_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1270_out;
SharedReg1311_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1311_out;
Delay102No8_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_3_cast <= Delay102No8_out;
SharedReg1263_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1263_out;
SharedReg1276_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1276_out;
SharedReg1288_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1288_out;
SharedReg21_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg21_out;
SharedReg1266_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1266_out;
SharedReg1017_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1017_out;
SharedReg1302_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1302_out;
Delay97No2_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_11_cast <= Delay97No2_out;
SharedReg320_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg320_out;
SharedReg1007_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1007_out;
   MUX_Product110_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1270_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1311_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay97No2_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg320_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1007_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay102No8_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1263_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1276_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1288_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg21_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1266_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1017_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1302_out_to_MUX_Product110_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_2_impl_1_out);

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_2_impl_1_out,
                 Y => Delay1No17_out);

Delay1No18_out_to_Product110_3_impl_parent_implementedSystem_port_0_cast <= Delay1No18_out;
Delay1No19_out_to_Product110_3_impl_parent_implementedSystem_port_1_cast <= Delay1No19_out;
   Product110_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_3_impl_out,
                 X => Delay1No18_out_to_Product110_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No19_out_to_Product110_3_impl_parent_implementedSystem_port_1_cast);

SharedReg856_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg856_out;
SharedReg429_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg429_out;
SharedReg1270_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1270_out;
SharedReg26_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg26_out;
SharedReg897_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg897_out;
Delay1No334_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_6_cast <= Delay1No334_out;
SharedReg384_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg384_out;
SharedReg794_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg794_out;
SharedReg791_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg791_out;
SharedReg379_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg379_out;
SharedReg1256_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1256_out;
SharedReg1302_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1302_out;
SharedReg654_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg654_out;
   MUX_Product110_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg856_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg429_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1256_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1302_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg654_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1270_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg26_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg897_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay1No334_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg384_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg794_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg791_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg379_out_to_MUX_Product110_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_3_impl_0_out);

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_3_impl_0_out,
                 Y => Delay1No18_out);

SharedReg1280_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1280_out;
SharedReg1098_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1098_out;
SharedReg1270_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1270_out;
SharedReg1003_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1003_out;
SharedReg1295_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1295_out;
SharedReg1263_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1263_out;
SharedReg1276_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1276_out;
SharedReg1288_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1288_out;
SharedReg32_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg32_out;
SharedReg1266_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1266_out;
SharedReg1127_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1127_out;
SharedReg1302_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1302_out;
Delay97No3_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_13_cast <= Delay97No3_out;
   MUX_Product110_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1280_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1098_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1127_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1302_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay97No3_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1270_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1003_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1295_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1263_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1276_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1288_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg32_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1266_out_to_MUX_Product110_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_3_impl_1_out);

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_3_impl_1_out,
                 Y => Delay1No19_out);

Delay1No20_out_to_Product110_4_impl_parent_implementedSystem_port_0_cast <= Delay1No20_out;
Delay1No21_out_to_Product110_4_impl_parent_implementedSystem_port_1_cast <= Delay1No21_out;
   Product110_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_4_impl_out,
                 X => Delay1No20_out_to_Product110_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No21_out_to_Product110_4_impl_parent_implementedSystem_port_1_cast);

SharedReg712_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg712_out;
SharedReg1317_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1317_out;
SharedReg1197_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1197_out;
SharedReg1094_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1094_out;
SharedReg100_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg100_out;
SharedReg1169_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1169_out;
SharedReg903_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg903_out;
Delay1No335_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_8_cast <= Delay1No335_out;
SharedReg393_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg393_out;
SharedReg855_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg855_out;
SharedReg800_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg800_out;
SharedReg386_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg386_out;
SharedReg1256_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1256_out;
   MUX_Product110_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg712_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1317_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg800_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg386_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1256_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1197_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1094_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg100_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1169_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg903_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay1No335_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg393_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg855_out_to_MUX_Product110_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_4_impl_0_out);

   Delay1No20_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_4_impl_0_out,
                 Y => Delay1No20_out);

Delay87No16_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_1_cast <= Delay87No16_out;
SharedReg1317_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1317_out;
SharedReg1280_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1280_out;
SharedReg1028_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1028_out;
SharedReg1029_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1029_out;
SharedReg1285_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1285_out;
SharedReg1295_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1295_out;
SharedReg1263_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1263_out;
SharedReg1276_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1276_out;
SharedReg1288_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1288_out;
SharedReg43_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg43_out;
SharedReg1266_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1266_out;
SharedReg965_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg965_out;
   MUX_Product110_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay87No16_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1317_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg43_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1266_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg965_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1280_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1028_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1029_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1285_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1295_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1263_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1276_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1288_out_to_MUX_Product110_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_4_impl_1_out);

   Delay1No21_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_4_impl_1_out,
                 Y => Delay1No21_out);

Delay1No22_out_to_Product110_5_impl_parent_implementedSystem_port_0_cast <= Delay1No22_out;
Delay1No23_out_to_Product110_5_impl_parent_implementedSystem_port_1_cast <= Delay1No23_out;
   Product110_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product110_5_impl_out,
                 X => Delay1No22_out_to_Product110_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No23_out_to_Product110_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1191_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1191_out;
SharedReg1315_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1315_out;
SharedReg1256_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1256_out;
SharedReg672_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg672_out;
SharedReg395_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg395_out;
SharedReg1181_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1181_out;
SharedReg907_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg907_out;
SharedReg449_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg449_out;
SharedReg50_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg50_out;
Delay1No342_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_10_cast <= Delay1No342_out;
SharedReg443_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg443_out;
SharedReg395_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg395_out;
SharedReg1194_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1194_out;
   MUX_Product110_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1191_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1315_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg443_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg395_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1194_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1256_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg672_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg395_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1181_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg907_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg449_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg50_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay1No342_out_to_MUX_Product110_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_5_impl_0_out);

   Delay1No22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_5_impl_0_out,
                 Y => Delay1No22_out);

SharedReg1266_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1266_out;
SharedReg1315_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1315_out;
SharedReg1115_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1115_out;
Delay87No17_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_4_cast <= Delay87No17_out;
SharedReg1294_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1294_out;
SharedReg1311_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1311_out;
SharedReg1284_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1284_out;
SharedReg1305_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1305_out;
SharedReg225_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg225_out;
SharedReg1263_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1263_out;
SharedReg1314_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1314_out;
SharedReg1288_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1288_out;
SharedReg1289_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1289_out;
   MUX_Product110_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1266_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1315_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1314_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1288_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1289_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1115_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay87No17_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1294_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1311_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1284_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1305_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg225_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1263_out_to_MUX_Product110_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product110_5_impl_1_out);

   Delay1No23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product110_5_impl_1_out,
                 Y => Delay1No23_out);

Delay1No24_out_to_Product109_0_impl_parent_implementedSystem_port_0_cast <= Delay1No24_out;
Delay1No25_out_to_Product109_0_impl_parent_implementedSystem_port_1_cast <= Delay1No25_out;
   Product109_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product109_0_impl_out,
                 X => Delay1No24_out_to_Product109_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No25_out_to_Product109_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1274_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1263_out;
SharedReg405_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg405_out;
SharedReg455_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg455_out;
SharedReg1256_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1256_out;
SharedReg1266_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1266_out;
SharedReg1267_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1267_out;
SharedReg1268_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1268_out;
SharedReg1269_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1269_out;
SharedReg727_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg727_out;
SharedReg1271_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1271_out;
SharedReg1299_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1299_out;
SharedReg1273_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1273_out;
   MUX_Product109_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1274_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1263_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1271_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1299_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1273_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg405_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg455_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1256_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1266_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1267_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1268_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1269_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg727_out_to_MUX_Product109_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_0_impl_0_out);

   Delay1No24_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_0_impl_0_out,
                 Y => Delay1No24_out);

SharedReg1274_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1263_out;
SharedReg1307_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1307_out;
SharedReg71_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg71_out;
SharedReg1139_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1139_out;
SharedReg1266_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1266_out;
SharedReg1267_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1267_out;
SharedReg1268_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1268_out;
SharedReg1269_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1269_out;
SharedReg1310_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1310_out;
SharedReg1271_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1271_out;
SharedReg1299_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1299_out;
SharedReg1273_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1273_out;
   MUX_Product109_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1274_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1263_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1271_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1299_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1273_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1307_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg71_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1139_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1266_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1267_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1268_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1269_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1310_out_to_MUX_Product109_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_0_impl_1_out);

   Delay1No25_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_0_impl_1_out,
                 Y => Delay1No25_out);

Delay1No26_out_to_Product109_1_impl_parent_implementedSystem_port_0_cast <= Delay1No26_out;
Delay1No27_out_to_Product109_1_impl_parent_implementedSystem_port_1_cast <= Delay1No27_out;
   Product109_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product109_1_impl_out,
                 X => Delay1No26_out_to_Product109_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No27_out_to_Product109_1_impl_parent_implementedSystem_port_1_cast);

SharedReg417_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg417_out;
SharedReg1305_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1305_out;
SharedReg1274_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1274_out;
SharedReg457_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg457_out;
SharedReg777_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg777_out;
SharedReg500_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg500_out;
SharedReg1256_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1256_out;
SharedReg1266_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1266_out;
SharedReg1267_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1267_out;
SharedReg1268_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1268_out;
SharedReg1269_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1269_out;
SharedReg786_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg786_out;
SharedReg1271_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1271_out;
   MUX_Product109_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg417_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1305_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1269_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg786_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1271_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1274_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg457_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg777_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg500_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1256_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1266_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1267_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1268_out_to_MUX_Product109_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_1_impl_0_out);

   Delay1No26_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_1_impl_0_out,
                 Y => Delay1No26_out);

Delay102No1_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_1_cast <= Delay102No1_out;
SharedReg1305_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1305_out;
SharedReg1274_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1274_out;
SharedReg1061_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1061_out;
SharedReg1289_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1289_out;
SharedReg194_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg194_out;
SharedReg1003_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1003_out;
SharedReg1266_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1266_out;
SharedReg1267_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1267_out;
SharedReg1268_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1268_out;
SharedReg1269_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1269_out;
SharedReg1310_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1310_out;
SharedReg1271_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1271_out;
   MUX_Product109_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay102No1_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1305_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1269_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1310_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1271_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1274_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1061_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1289_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg194_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1003_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1266_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1267_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1268_out_to_MUX_Product109_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_1_impl_1_out);

   Delay1No27_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_1_impl_1_out,
                 Y => Delay1No27_out);

Delay1No28_out_to_Product109_2_impl_parent_implementedSystem_port_0_cast <= Delay1No28_out;
Delay1No29_out_to_Product109_2_impl_parent_implementedSystem_port_1_cast <= Delay1No29_out;
   Product109_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product109_2_impl_out,
                 X => Delay1No28_out_to_Product109_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No29_out_to_Product109_2_impl_parent_implementedSystem_port_1_cast);

SharedReg797_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg797_out;
SharedReg508_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg508_out;
Delay87No8_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_3_cast <= Delay87No8_out;
SharedReg1273_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1273_out;
SharedReg888_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg888_out;
SharedReg836_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg836_out;
SharedReg784_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg784_out;
SharedReg505_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg505_out;
SharedReg1256_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1256_out;
SharedReg1266_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1266_out;
SharedReg1267_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1267_out;
SharedReg1268_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1268_out;
SharedReg1269_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1269_out;
   MUX_Product109_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg797_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg508_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1267_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1268_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1269_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay87No8_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1273_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg888_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg836_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg784_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg505_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1256_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1266_out_to_MUX_Product109_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_2_impl_0_out);

   Delay1No28_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_2_impl_0_out,
                 Y => Delay1No28_out);

SharedReg1294_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1294_out;
SharedReg1271_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1271_out;
Delay102No2_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_3_cast <= Delay102No2_out;
SharedReg1273_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1273_out;
SharedReg1314_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1314_out;
SharedReg1288_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1288_out;
SharedReg1289_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1289_out;
SharedReg205_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg205_out;
SharedReg1129_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1129_out;
SharedReg1266_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1266_out;
SharedReg1267_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1267_out;
SharedReg1268_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1268_out;
SharedReg1269_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1269_out;
   MUX_Product109_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1294_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1271_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1267_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1268_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1269_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay102No2_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1273_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1314_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1288_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1289_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg205_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1129_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1266_out_to_MUX_Product109_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_2_impl_1_out);

   Delay1No29_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_2_impl_1_out,
                 Y => Delay1No29_out);

Delay1No30_out_to_Product109_3_impl_parent_implementedSystem_port_0_cast <= Delay1No30_out;
Delay1No31_out_to_Product109_3_impl_parent_implementedSystem_port_1_cast <= Delay1No31_out;
   Product109_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product109_3_impl_out,
                 X => Delay1No30_out_to_Product109_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No31_out_to_Product109_3_impl_parent_implementedSystem_port_1_cast);

SharedReg653_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg653_out;
SharedReg803_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg803_out;
SharedReg805_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg805_out;
SharedReg801_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg801_out;
SharedReg28_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg28_out;
Delay1No340_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_6_cast <= Delay1No340_out;
SharedReg1161_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1161_out;
SharedReg895_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg895_out;
SharedReg845_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg845_out;
SharedReg653_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg653_out;
SharedReg1256_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1256_out;
SharedReg1266_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1266_out;
SharedReg1267_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1267_out;
   MUX_Product109_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg653_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg803_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1256_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1266_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1267_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg805_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg801_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg28_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay1No340_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1161_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg895_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg845_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg653_out_to_MUX_Product109_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_3_impl_0_out);

   Delay1No30_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_3_impl_0_out,
                 Y => Delay1No30_out);

SharedReg329_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg329_out;
SharedReg1098_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1098_out;
SharedReg1294_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1294_out;
SharedReg1311_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1311_out;
SharedReg203_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg203_out;
SharedReg1263_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1263_out;
SharedReg1314_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1314_out;
SharedReg1288_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1288_out;
SharedReg1289_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1289_out;
SharedReg216_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg216_out;
SharedReg967_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg967_out;
SharedReg1266_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1266_out;
SharedReg1267_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1267_out;
   MUX_Product109_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg329_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1098_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg967_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1266_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1267_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1294_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1311_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg203_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1263_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1314_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1288_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1289_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg216_out_to_MUX_Product109_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_3_impl_1_out);

   Delay1No31_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_3_impl_1_out,
                 Y => Delay1No31_out);

Delay1No32_out_to_Product109_4_impl_parent_implementedSystem_port_0_cast <= Delay1No32_out;
Delay1No33_out_to_Product109_4_impl_parent_implementedSystem_port_1_cast <= Delay1No33_out;
   Product109_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product109_4_impl_out,
                 X => Delay1No32_out_to_Product109_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No33_out_to_Product109_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1302_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1302_out;
SharedReg663_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg663_out;
SharedReg662_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg662_out;
SharedReg570_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg570_out;
SharedReg901_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg901_out;
SharedReg441_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg441_out;
SharedReg39_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg39_out;
Delay1No341_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_8_cast <= Delay1No341_out;
SharedReg387_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg387_out;
SharedReg1169_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1169_out;
SharedReg902_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg902_out;
SharedReg662_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg662_out;
SharedReg1256_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1256_out;
   MUX_Product109_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1302_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg663_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg902_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg662_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1256_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg662_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg570_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg901_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg441_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg39_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay1No341_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg387_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1169_out_to_MUX_Product109_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_4_impl_0_out);

   Delay1No32_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_4_impl_0_out,
                 Y => Delay1No32_out);

SharedReg1302_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1302_out;
Delay97No4_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_2_cast <= Delay97No4_out;
SharedReg338_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg338_out;
SharedReg973_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg973_out;
SharedReg1284_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1284_out;
SharedReg1305_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1305_out;
SharedReg214_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg214_out;
SharedReg1263_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1263_out;
SharedReg1314_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1314_out;
SharedReg1288_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1288_out;
SharedReg1289_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1289_out;
SharedReg227_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg227_out;
SharedReg969_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg969_out;
   MUX_Product109_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1302_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay97No4_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1289_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg227_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg969_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg338_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg973_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1284_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1305_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg214_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1263_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1314_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1288_out_to_MUX_Product109_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_4_impl_1_out);

   Delay1No33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_4_impl_1_out,
                 Y => Delay1No33_out);

Delay1No34_out_to_Product109_5_impl_parent_implementedSystem_port_0_cast <= Delay1No34_out;
Delay1No35_out_to_Product109_5_impl_parent_implementedSystem_port_1_cast <= Delay1No35_out;
   Product109_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product109_5_impl_out,
                 X => Delay1No34_out_to_Product109_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No35_out_to_Product109_5_impl_parent_implementedSystem_port_1_cast);

SharedReg56_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg56_out;
SharedReg625_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg625_out;
SharedReg1256_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1256_out;
SharedReg1302_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1302_out;
SharedReg281_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg281_out;
SharedReg968_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg968_out;
SharedReg908_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg908_out;
SharedReg48_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg48_out;
SharedReg1192_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1192_out;
Delay1No348_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_10_cast <= Delay1No348_out;
SharedReg1273_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1273_out;
SharedReg1306_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1306_out;
SharedReg1300_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1300_out;
   MUX_Product109_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg56_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg625_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1273_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1306_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1300_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1256_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1302_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg281_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg968_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg908_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg48_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1192_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay1No348_out_to_MUX_Product109_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_5_impl_0_out);

   Delay1No34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_5_impl_0_out,
                 Y => Delay1No34_out);

SharedReg230_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg230_out;
SharedReg121_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg121_out;
SharedReg1046_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1046_out;
SharedReg1302_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1302_out;
SharedReg221_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg221_out;
SharedReg1115_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1115_out;
SharedReg1272_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1272_out;
SharedReg969_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg969_out;
SharedReg1274_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1263_out;
SharedReg1273_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1273_out;
SharedReg1306_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1306_out;
SharedReg1300_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1300_out;
   MUX_Product109_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg230_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg121_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1273_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1306_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1300_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1046_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1302_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg221_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1115_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1272_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg969_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1274_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1263_out_to_MUX_Product109_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product109_5_impl_1_out);

   Delay1No35_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product109_5_impl_1_out,
                 Y => Delay1No35_out);

Delay1No36_out_to_Product111_0_impl_parent_implementedSystem_port_0_cast <= Delay1No36_out;
Delay1No37_out_to_Product111_0_impl_parent_implementedSystem_port_1_cast <= Delay1No37_out;
   Product111_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_0_impl_out,
                 X => Delay1No36_out_to_Product111_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No37_out_to_Product111_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1313_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1313_out;
SharedReg1263_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1263_out;
SharedReg1264_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1264_out;
SharedReg450_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg450_out;
SharedReg1256_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1256_out;
SharedReg1308_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1308_out;
SharedReg679_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg679_out;
Delay62No_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_8_cast <= Delay62No_out;
SharedReg537_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg537_out;
SharedReg1282_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1282_out;
SharedReg1137_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1137_out;
SharedReg1312_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1312_out;
SharedReg531_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg531_out;
   MUX_Product111_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1313_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1263_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1137_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1312_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg531_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1264_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg450_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1256_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1308_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg679_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay62No_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg537_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1282_out_to_MUX_Product111_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_0_impl_0_out);

   Delay1No36_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_0_impl_0_out,
                 Y => Delay1No36_out);

SharedReg1313_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1313_out;
SharedReg1263_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1263_out;
SharedReg1264_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1264_out;
SharedReg305_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg305_out;
SharedReg1082_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1082_out;
SharedReg1308_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1308_out;
SharedReg1317_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1317_out;
SharedReg9_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg9_out;
SharedReg1088_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1088_out;
SharedReg1282_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1282_out;
SharedReg977_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg977_out;
SharedReg1312_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1312_out;
SharedReg1089_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1089_out;
   MUX_Product111_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1313_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1263_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg977_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1312_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1089_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1264_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg305_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1082_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1308_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1317_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg9_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1088_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1282_out_to_MUX_Product111_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_0_impl_1_out);

   Delay1No37_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_0_impl_1_out,
                 Y => Delay1No37_out);

Delay1No38_out_to_Product111_1_impl_parent_implementedSystem_port_0_cast <= Delay1No38_out;
Delay1No39_out_to_Product111_1_impl_parent_implementedSystem_port_1_cast <= Delay1No39_out;
   Product111_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_1_impl_out,
                 X => Delay1No38_out_to_Product111_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No39_out_to_Product111_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1299_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1299_out;
SharedReg1273_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1273_out;
SharedReg1313_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1313_out;
SharedReg1263_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1263_out;
SharedReg12_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg12_out;
SharedReg1315_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1315_out;
SharedReg1256_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1256_out;
SharedReg1308_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1308_out;
SharedReg737_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg737_out;
SharedReg462_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg462_out;
SharedReg546_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg546_out;
SharedReg1282_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1282_out;
SharedReg1059_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1059_out;
   MUX_Product111_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1299_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1273_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg546_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1282_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1059_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1313_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1263_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg12_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1315_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1256_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1308_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg737_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg462_out_to_MUX_Product111_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_1_impl_0_out);

   Delay1No38_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_1_impl_0_out,
                 Y => Delay1No38_out);

SharedReg1299_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1299_out;
SharedReg1273_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1273_out;
SharedReg1313_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1313_out;
SharedReg1263_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1263_out;
SharedReg186_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg186_out;
SharedReg1315_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1315_out;
SharedReg933_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg933_out;
SharedReg1308_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1308_out;
SharedReg1317_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1317_out;
SharedReg20_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg20_out;
SharedReg939_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg939_out;
SharedReg1282_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1282_out;
SharedReg991_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg991_out;
   MUX_Product111_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1299_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1273_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg939_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1282_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg991_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1313_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1263_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg186_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1315_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg933_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1308_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1317_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg20_out_to_MUX_Product111_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_1_impl_1_out);

   Delay1No39_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_1_impl_1_out,
                 Y => Delay1No39_out);

Delay1No40_out_to_Product111_2_impl_parent_implementedSystem_port_0_cast <= Delay1No40_out;
Delay1No41_out_to_Product111_2_impl_parent_implementedSystem_port_1_cast <= Delay1No41_out;
   Product111_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_2_impl_out,
                 X => Delay1No40_out_to_Product111_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No41_out_to_Product111_2_impl_parent_implementedSystem_port_1_cast);

SharedReg846_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg846_out;
SharedReg1271_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1271_out;
SharedReg1299_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1299_out;
SharedReg1305_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1305_out;
SharedReg1306_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1306_out;
SharedReg1300_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1300_out;
SharedReg23_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg23_out;
SharedReg1315_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1315_out;
SharedReg1256_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1256_out;
SharedReg1308_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1308_out;
SharedReg750_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg750_out;
SharedReg467_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg467_out;
SharedReg555_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg555_out;
   MUX_Product111_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg846_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1271_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg750_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg467_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg555_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1299_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1305_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1306_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1300_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg23_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1315_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1256_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1308_out_to_MUX_Product111_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_2_impl_0_out);

   Delay1No40_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_2_impl_0_out,
                 Y => Delay1No40_out);

SharedReg1310_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1310_out;
SharedReg1271_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1271_out;
SharedReg1299_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1299_out;
SharedReg1305_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1305_out;
SharedReg1306_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1306_out;
SharedReg1300_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1300_out;
SharedReg197_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg197_out;
SharedReg1315_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1315_out;
SharedReg943_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg943_out;
SharedReg1308_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1308_out;
SharedReg1317_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1317_out;
SharedReg31_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg31_out;
SharedReg949_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg949_out;
   MUX_Product111_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1310_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1271_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1317_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg31_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg949_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1299_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1305_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1306_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1300_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg197_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1315_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg943_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1308_out_to_MUX_Product111_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_2_impl_1_out);

   Delay1No41_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_2_impl_1_out,
                 Y => Delay1No41_out);

Delay1No42_out_to_Product111_3_impl_parent_implementedSystem_port_0_cast <= Delay1No42_out;
Delay1No43_out_to_Product111_3_impl_parent_implementedSystem_port_1_cast <= Delay1No43_out;
   Product111_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_3_impl_out,
                 X => Delay1No42_out_to_Product111_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No43_out_to_Product111_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1268_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1268_out;
SharedReg1269_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1269_out;
SharedReg1172_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1172_out;
SharedReg514_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg514_out;
SharedReg894_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg894_out;
Delay1No346_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_6_cast <= Delay1No346_out;
SharedReg1306_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1306_out;
SharedReg1300_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1300_out;
SharedReg34_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg34_out;
SharedReg1315_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1315_out;
SharedReg1256_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1256_out;
SharedReg1308_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1308_out;
SharedReg903_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg903_out;
   MUX_Product111_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1268_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1269_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1256_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1308_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg903_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1172_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg514_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg894_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay1No346_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1306_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1300_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg34_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1315_out_to_MUX_Product111_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_3_impl_0_out);

   Delay1No42_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_3_impl_0_out,
                 Y => Delay1No42_out);

SharedReg1268_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1268_out;
SharedReg1269_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1269_out;
SharedReg1310_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1310_out;
SharedReg1271_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1271_out;
SharedReg1274_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1263_out;
SharedReg1306_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1306_out;
SharedReg1300_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1300_out;
SharedReg208_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg208_out;
SharedReg1315_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1315_out;
SharedReg1091_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1091_out;
SharedReg1308_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1308_out;
SharedReg1317_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1317_out;
   MUX_Product111_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1268_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1269_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1091_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1308_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1317_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1310_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1271_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1274_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1263_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1306_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1300_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg208_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1315_out_to_MUX_Product111_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_3_impl_1_out);

   Delay1No43_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_3_impl_1_out,
                 Y => Delay1No43_out);

Delay1No44_out_to_Product111_4_impl_parent_implementedSystem_port_0_cast <= Delay1No44_out;
Delay1No45_out_to_Product111_4_impl_parent_implementedSystem_port_1_cast <= Delay1No45_out;
   Product111_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_4_impl_out,
                 X => Delay1No44_out_to_Product111_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No45_out_to_Product111_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1266_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1266_out;
SharedReg1267_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1267_out;
SharedReg1268_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1268_out;
SharedReg813_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg813_out;
SharedReg853_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg853_out;
SharedReg37_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg37_out;
SharedReg1168_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1168_out;
Delay1No347_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_8_cast <= Delay1No347_out;
SharedReg1306_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1306_out;
SharedReg1300_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1300_out;
SharedReg45_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg45_out;
SharedReg1315_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1315_out;
SharedReg1256_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1256_out;
   MUX_Product111_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1266_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1267_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg45_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1315_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1256_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1268_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg813_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg853_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg37_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1168_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay1No347_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1306_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1300_out_to_MUX_Product111_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_4_impl_0_out);

   Delay1No44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_4_impl_0_out,
                 Y => Delay1No44_out);

SharedReg1266_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1266_out;
SharedReg1267_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1267_out;
SharedReg1268_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1268_out;
SharedReg973_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg973_out;
SharedReg1272_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1272_out;
SharedReg1095_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1095_out;
SharedReg1274_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1263_out;
SharedReg1306_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1306_out;
SharedReg1300_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1300_out;
SharedReg219_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg219_out;
SharedReg1315_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1315_out;
SharedReg1094_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1094_out;
   MUX_Product111_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1266_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1267_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg219_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1315_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1094_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1268_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg973_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1272_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1095_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1274_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1263_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1306_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1300_out_to_MUX_Product111_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_4_impl_1_out);

   Delay1No45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_4_impl_1_out,
                 Y => Delay1No45_out);

Delay1No46_out_to_Product111_5_impl_parent_implementedSystem_port_0_cast <= Delay1No46_out;
Delay1No47_out_to_Product111_5_impl_parent_implementedSystem_port_1_cast <= Delay1No47_out;
   Product111_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product111_5_impl_out,
                 X => Delay1No46_out_to_Product111_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No47_out_to_Product111_5_impl_parent_implementedSystem_port_1_cast);

SharedReg117_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg117_out;
SharedReg573_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg573_out;
SharedReg1256_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1256_out;
SharedReg1266_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1266_out;
SharedReg1317_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1317_out;
SharedReg1187_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1187_out;
SharedReg527_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg527_out;
SharedReg1270_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1270_out;
SharedReg872_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg872_out;
SharedReg525_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg525_out;
SharedReg1305_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1305_out;
SharedReg1274_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1274_out;
SharedReg620_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg620_out;
   MUX_Product111_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg117_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg573_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1305_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1274_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg620_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1256_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1266_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1317_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1187_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg527_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1270_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg872_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg525_out_to_MUX_Product111_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_5_impl_0_out);

   Delay1No46_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_5_impl_0_out,
                 Y => Delay1No46_out);

SharedReg167_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg167_out;
SharedReg350_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg350_out;
SharedReg1070_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1070_out;
SharedReg1266_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1266_out;
SharedReg1317_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1317_out;
SharedReg1280_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1280_out;
SharedReg1251_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1251_out;
SharedReg1270_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1270_out;
SharedReg1311_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1311_out;
Delay102No11_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_10_cast <= Delay102No11_out;
SharedReg1305_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1305_out;
SharedReg1274_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1274_out;
SharedReg1107_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1107_out;
   MUX_Product111_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg167_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg350_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1305_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1274_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1107_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1070_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1266_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1317_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1280_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1251_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1270_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1311_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay102No11_out_to_MUX_Product111_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product111_5_impl_1_out);

   Delay1No47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product111_5_impl_1_out,
                 Y => Delay1No47_out);

Delay1No48_out_to_Product210_0_impl_parent_implementedSystem_port_0_cast <= Delay1No48_out;
Delay1No49_out_to_Product210_0_impl_parent_implementedSystem_port_1_cast <= Delay1No49_out;
   Product210_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_0_impl_out,
                 X => Delay1No48_out_to_Product210_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No49_out_to_Product210_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1274_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1263_out;
SharedReg495_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg495_out;
SharedReg1265_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1265_out;
SharedReg1256_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1256_out;
SharedReg1266_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1266_out;
SharedReg453_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg453_out;
SharedReg357_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg357_out;
SharedReg1293_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1293_out;
SharedReg400_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg400_out;
SharedReg1082_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1082_out;
SharedReg1272_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1272_out;
SharedReg539_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg539_out;
   MUX_Product210_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1274_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1263_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1082_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1272_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg539_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg495_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1265_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1256_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1266_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg453_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg357_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1293_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg400_out_to_MUX_Product210_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_0_impl_0_out);

   Delay1No48_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_0_impl_0_out,
                 Y => Delay1No48_out);

SharedReg1274_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1263_out;
SharedReg308_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg308_out;
SharedReg1265_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1265_out;
SharedReg940_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg940_out;
SharedReg1266_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1266_out;
SharedReg306_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg306_out;
SharedReg73_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg73_out;
SharedReg1293_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1293_out;
SharedReg1144_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1144_out;
SharedReg303_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg303_out;
SharedReg1272_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1272_out;
SharedReg984_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg984_out;
   MUX_Product210_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1274_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1263_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg303_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1272_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg984_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg308_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1265_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg940_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1266_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg306_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg73_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1293_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1144_out_to_MUX_Product210_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_0_impl_1_out);

   Delay1No49_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_0_impl_1_out,
                 Y => Delay1No49_out);

Delay1No50_out_to_Product210_1_impl_parent_implementedSystem_port_0_cast <= Delay1No50_out;
Delay1No51_out_to_Product210_1_impl_parent_implementedSystem_port_1_cast <= Delay1No51_out;
   Product210_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_1_impl_out,
                 X => Delay1No50_out_to_Product210_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No51_out_to_Product210_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1312_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1312_out;
SharedReg540_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg540_out;
SharedReg1274_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1263_out;
SharedReg77_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg77_out;
SharedReg461_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg461_out;
SharedReg1256_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1256_out;
SharedReg1266_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1266_out;
SharedReg458_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg458_out;
SharedReg366_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg366_out;
SharedReg1293_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1293_out;
SharedReg408_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg408_out;
SharedReg933_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg933_out;
   MUX_Product210_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1312_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg540_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1293_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg408_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg933_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1274_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1263_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg77_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg461_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1256_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1266_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg458_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg366_out_to_MUX_Product210_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_1_impl_0_out);

   Delay1No50_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_1_impl_0_out,
                 Y => Delay1No50_out);

SharedReg1312_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1312_out;
SharedReg941_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg941_out;
SharedReg1274_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1263_out;
SharedReg135_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg135_out;
SharedReg81_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg81_out;
SharedReg951_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg951_out;
SharedReg1266_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1266_out;
SharedReg315_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg315_out;
SharedReg83_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg83_out;
SharedReg1293_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1293_out;
SharedReg1066_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1066_out;
SharedReg312_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg312_out;
   MUX_Product210_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1312_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg941_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1293_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1066_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg312_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1274_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1263_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg135_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg81_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg951_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1266_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg315_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg83_out_to_MUX_Product210_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_1_impl_1_out);

   Delay1No51_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_1_impl_1_out,
                 Y => Delay1No51_out);

Delay1No52_out_to_Product210_2_impl_parent_implementedSystem_port_0_cast <= Delay1No52_out;
Delay1No53_out_to_Product210_2_impl_parent_implementedSystem_port_1_cast <= Delay1No53_out;
   Product210_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_2_impl_out,
                 X => Delay1No52_out_to_Product210_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No53_out_to_Product210_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1282_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1282_out;
SharedReg1017_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1017_out;
SharedReg1312_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1312_out;
SharedReg1273_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1273_out;
SharedReg1274_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1274_out;
SharedReg464_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg464_out;
SharedReg87_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg87_out;
SharedReg466_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg466_out;
SharedReg1256_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1256_out;
SharedReg1266_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1266_out;
SharedReg509_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg509_out;
SharedReg507_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg507_out;
SharedReg1293_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1293_out;
   MUX_Product210_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1282_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1017_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg509_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg507_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1293_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1312_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1273_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1274_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg464_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg87_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg466_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1256_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1266_out_to_MUX_Product210_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_2_impl_0_out);

   Delay1No52_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_2_impl_0_out,
                 Y => Delay1No52_out);

SharedReg1282_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1282_out;
SharedReg1002_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1002_out;
SharedReg1312_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1312_out;
SharedReg1273_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1273_out;
SharedReg1274_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1274_out;
SharedReg1020_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1020_out;
SharedReg143_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg143_out;
SharedReg91_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg91_out;
SharedReg961_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg961_out;
SharedReg1266_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1266_out;
SharedReg324_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg324_out;
SharedReg93_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg93_out;
SharedReg1293_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1293_out;
   MUX_Product210_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1282_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1002_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg324_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg93_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1293_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1312_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1273_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1274_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1020_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg143_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg91_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg961_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1266_out_to_MUX_Product210_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_2_impl_1_out);

   Delay1No53_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_2_impl_1_out,
                 Y => Delay1No53_out);

Delay1No54_out_to_Product210_3_impl_parent_implementedSystem_port_0_cast <= Delay1No54_out;
Delay1No55_out_to_Product210_3_impl_parent_implementedSystem_port_1_cast <= Delay1No55_out;
   Product210_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_3_impl_out,
                 X => Delay1No54_out_to_Product210_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No55_out_to_Product210_3_impl_parent_implementedSystem_port_1_cast);

SharedReg516_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg516_out;
SharedReg562_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg562_out;
SharedReg1282_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1282_out;
SharedReg1271_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1271_out;
SharedReg380_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg380_out;
SharedReg1273_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1273_out;
SharedReg1274_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1274_out;
SharedReg512_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg512_out;
SharedReg97_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg97_out;
SharedReg475_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg475_out;
SharedReg1256_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1256_out;
SharedReg1266_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1266_out;
SharedReg560_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg560_out;
   MUX_Product210_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg516_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg562_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1256_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1266_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg560_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1282_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1271_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg380_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1273_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1274_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg512_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg97_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg475_out_to_MUX_Product210_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_3_impl_0_out);

   Delay1No54_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_3_impl_0_out,
                 Y => Delay1No54_out);

SharedReg42_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg42_out;
SharedReg1134_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1134_out;
SharedReg1282_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1282_out;
SharedReg1271_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1271_out;
Delay102No9_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_5_cast <= Delay102No9_out;
SharedReg1273_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1273_out;
SharedReg1274_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1274_out;
SharedReg1031_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1031_out;
SharedReg151_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg151_out;
SharedReg101_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg101_out;
SharedReg1100_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1100_out;
SharedReg1266_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1266_out;
SharedReg333_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg333_out;
   MUX_Product210_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg42_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1134_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1100_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1266_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg333_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1282_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1271_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay102No9_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1273_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1274_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1031_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg151_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg101_out_to_MUX_Product210_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_3_impl_1_out);

   Delay1No55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_3_impl_1_out,
                 Y => Delay1No55_out);

Delay1No56_out_to_Product210_4_impl_parent_implementedSystem_port_0_cast <= Delay1No56_out;
Delay1No57_out_to_Product210_4_impl_parent_implementedSystem_port_1_cast <= Delay1No57_out;
   Product210_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_4_impl_out,
                 X => Delay1No56_out_to_Product210_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No57_out_to_Product210_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1308_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1308_out;
SharedReg910_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg910_out;
SharedReg523_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg523_out;
SharedReg1269_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1269_out;
SharedReg1270_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1270_out;
SharedReg863_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg863_out;
SharedReg434_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg434_out;
SharedReg1273_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1273_out;
SharedReg1274_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1274_out;
SharedReg568_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg568_out;
SharedReg107_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg107_out;
SharedReg521_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg521_out;
SharedReg1256_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1256_out;
   MUX_Product210_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1308_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg910_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg107_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg521_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1256_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg523_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1269_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1270_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg863_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg434_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1273_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1274_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg568_out_to_MUX_Product210_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_4_impl_0_out);

   Delay1No56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_4_impl_0_out,
                 Y => Delay1No56_out);

SharedReg1308_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1308_out;
SharedReg1317_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1317_out;
SharedReg53_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg53_out;
SharedReg1269_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1269_out;
SharedReg1270_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1270_out;
SharedReg1311_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1311_out;
Delay102No10_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_7_cast <= Delay102No10_out;
SharedReg1273_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1273_out;
SharedReg1274_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1274_out;
SharedReg1118_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1118_out;
SharedReg159_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg159_out;
SharedReg111_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg111_out;
SharedReg1077_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1077_out;
   MUX_Product210_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1308_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1317_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg159_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg111_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1077_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg53_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1269_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1270_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1311_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay102No10_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1273_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1274_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1118_out_to_MUX_Product210_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_4_impl_1_out);

   Delay1No57_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_4_impl_1_out,
                 Y => Delay1No57_out);

Delay1No58_out_to_Product210_5_impl_parent_implementedSystem_port_0_cast <= Delay1No58_out;
Delay1No59_out_to_Product210_5_impl_parent_implementedSystem_port_1_cast <= Delay1No59_out;
   Product210_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product210_5_impl_out,
                 X => Delay1No58_out_to_Product210_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No59_out_to_Product210_5_impl_parent_implementedSystem_port_1_cast);

SharedReg529_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg529_out;
SharedReg1265_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1265_out;
SharedReg1256_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1256_out;
SharedReg1308_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1308_out;
SharedReg620_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg620_out;
SharedReg619_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg619_out;
SharedReg774_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg774_out;
SharedReg725_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg725_out;
SharedReg491_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg491_out;
Delay87No11_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_10_cast <= Delay87No11_out;
SharedReg1273_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1273_out;
SharedReg1274_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1263_out;
   MUX_Product210_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg529_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1265_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1273_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1274_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1263_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1256_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1308_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg620_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg619_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg774_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg725_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg491_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay87No11_out_to_MUX_Product210_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_5_impl_0_out);

   Delay1No58_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_5_impl_0_out,
                 Y => Delay1No58_out);

SharedReg1307_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1307_out;
SharedReg1265_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1265_out;
SharedReg1052_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1052_out;
SharedReg1308_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1308_out;
Delay97No5_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_5_cast <= Delay97No5_out;
SharedReg347_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg347_out;
SharedReg1251_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1251_out;
SharedReg1294_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1294_out;
SharedReg1271_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1271_out;
Delay102No5_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_10_cast <= Delay102No5_out;
SharedReg1273_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1273_out;
SharedReg1274_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1263_out;
   MUX_Product210_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1307_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1265_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1273_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1274_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1263_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1052_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1308_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay97No5_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg347_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1251_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1294_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1271_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay102No5_out_to_MUX_Product210_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product210_5_impl_1_out);

   Delay1No59_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product210_5_impl_1_out,
                 Y => Delay1No59_out);

Delay1No60_out_to_Product310_0_impl_parent_implementedSystem_port_0_cast <= Delay1No60_out;
Delay1No61_out_to_Product310_0_impl_parent_implementedSystem_port_1_cast <= Delay1No61_out;
   Product310_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_0_impl_out,
                 X => Delay1No60_out_to_Product310_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No61_out_to_Product310_0_impl_parent_implementedSystem_port_1_cast);

SharedReg536_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg536_out;
SharedReg493_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg493_out;
SharedReg531_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg531_out;
SharedReg680_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg680_out;
SharedReg1256_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1256_out;
SharedReg402_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg402_out;
SharedReg497_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg497_out;
SharedReg400_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg400_out;
SharedReg538_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg538_out;
SharedReg450_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg450_out;
SharedReg1082_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1082_out;
SharedReg1272_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1272_out;
SharedReg130_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg130_out;
   MUX_Product310_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg536_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg493_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1082_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1272_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg130_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg531_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg680_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1256_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg402_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg497_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg400_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg538_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg450_out_to_MUX_Product310_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_0_impl_0_out);

   Delay1No60_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_0_impl_0_out,
                 Y => Delay1No60_out);

SharedReg132_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg132_out;
SharedReg1275_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1275_out;
SharedReg179_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg179_out;
Delay94No_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_4_cast <= Delay94No_out;
SharedReg1059_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1059_out;
SharedReg1146_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1146_out;
SharedReg1087_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1087_out;
SharedReg75_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg75_out;
SharedReg1142_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1142_out;
SharedReg129_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg129_out;
SharedReg977_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg977_out;
SharedReg1272_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1272_out;
SharedReg978_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg978_out;
   MUX_Product310_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg132_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1275_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg977_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1272_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg978_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg179_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay94No_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1059_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1146_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1087_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg75_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1142_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg129_out_to_MUX_Product310_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_0_impl_1_out);

   Delay1No61_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_0_impl_1_out,
                 Y => Delay1No61_out);

Delay1No62_out_to_Product310_1_impl_parent_implementedSystem_port_0_cast <= Delay1No62_out;
Delay1No63_out_to_Product310_1_impl_parent_implementedSystem_port_1_cast <= Delay1No63_out;
   Product310_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_1_impl_out,
                 X => Delay1No62_out_to_Product310_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No63_out_to_Product310_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1272_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1272_out;
Delay19No7_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_2_cast <= Delay19No7_out;
SharedReg545_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg545_out;
SharedReg1263_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1263_out;
SharedReg549_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg549_out;
SharedReg499_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg499_out;
SharedReg1256_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1256_out;
SharedReg457_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg457_out;
SharedReg547_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg547_out;
SharedReg499_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg499_out;
SharedReg596_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg596_out;
SharedReg456_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg456_out;
SharedReg933_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg933_out;
   MUX_Product310_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1272_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay19No7_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg596_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg456_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg933_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg545_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1263_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg549_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg499_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1256_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg457_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg547_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg499_out_to_MUX_Product310_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_1_impl_0_out);

   Delay1No62_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_1_impl_0_out,
                 Y => Delay1No62_out);

SharedReg1272_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1272_out;
SharedReg997_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg997_out;
SharedReg140_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg140_out;
SharedReg1263_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1263_out;
SharedReg1307_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1307_out;
SharedReg314_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg314_out;
SharedReg1017_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1017_out;
SharedReg1069_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1069_out;
SharedReg938_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg938_out;
SharedReg85_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg85_out;
SharedReg1064_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1064_out;
SharedReg137_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg137_out;
SharedReg991_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg991_out;
   MUX_Product310_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1272_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg997_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1064_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg137_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg991_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg140_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1263_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1307_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg314_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1017_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1069_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg938_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg85_out_to_MUX_Product310_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_1_impl_1_out);

   Delay1No63_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_1_impl_1_out,
                 Y => Delay1No63_out);

Delay1No64_out_to_Product310_2_impl_parent_implementedSystem_port_0_cast <= Delay1No64_out;
Delay1No65_out_to_Product310_2_impl_parent_implementedSystem_port_1_cast <= Delay1No65_out;
   Product310_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_2_impl_out,
                 X => Delay1No64_out_to_Product310_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No65_out_to_Product310_2_impl_parent_implementedSystem_port_1_cast);

SharedReg418_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg418_out;
SharedReg943_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg943_out;
SharedReg1272_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1272_out;
SharedReg550_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg550_out;
SharedReg1274_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1263_out;
SharedReg556_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg556_out;
SharedReg550_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg550_out;
SharedReg1256_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1256_out;
SharedReg506_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg506_out;
SharedReg650_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg650_out;
SharedReg504_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg504_out;
SharedReg698_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg698_out;
   MUX_Product310_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg418_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg943_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg650_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg504_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg698_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1272_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg550_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1274_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1263_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg556_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg550_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1256_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg506_out_to_MUX_Product310_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_2_impl_0_out);

   Delay1No64_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_2_impl_0_out,
                 Y => Delay1No64_out);

SharedReg1025_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1025_out;
SharedReg321_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg321_out;
SharedReg1272_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1272_out;
SharedReg952_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg952_out;
SharedReg1274_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1263_out;
SharedReg1307_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1307_out;
SharedReg323_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg323_out;
SharedReg1091_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1091_out;
SharedReg1027_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1027_out;
SharedReg948_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg948_out;
SharedReg95_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg95_out;
SharedReg1023_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1023_out;
   MUX_Product310_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1025_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg321_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg948_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg95_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1023_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1272_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg952_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1274_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1263_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1307_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg323_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1091_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1027_out_to_MUX_Product310_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_2_impl_1_out);

   Delay1No65_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_2_impl_1_out,
                 Y => Delay1No65_out);

Delay1No66_out_to_Product310_3_impl_parent_implementedSystem_port_0_cast <= Delay1No66_out;
Delay1No67_out_to_Product310_3_impl_parent_implementedSystem_port_1_cast <= Delay1No67_out;
   Product310_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_3_impl_out,
                 X => Delay1No66_out_to_Product310_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No67_out_to_Product310_3_impl_parent_implementedSystem_port_1_cast);

SharedReg513_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg513_out;
SharedReg1293_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1293_out;
SharedReg425_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg425_out;
SharedReg1028_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1028_out;
Delay87No9_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_5_cast <= Delay87No9_out;
SharedReg1305_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1305_out;
SharedReg1274_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1263_out;
SharedReg564_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg564_out;
SharedReg652_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg652_out;
SharedReg1256_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1256_out;
SharedReg607_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg607_out;
SharedReg659_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg659_out;
   MUX_Product310_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg513_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1293_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1256_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg607_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg659_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg425_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1028_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay87No9_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1305_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1274_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1263_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg564_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg652_out_to_MUX_Product310_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_3_impl_0_out);

   Delay1No66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_3_impl_0_out,
                 Y => Delay1No66_out);

SharedReg103_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg103_out;
SharedReg1293_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1293_out;
SharedReg1039_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1039_out;
SharedReg1094_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1094_out;
Delay102No3_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_5_cast <= Delay102No3_out;
SharedReg1305_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1305_out;
SharedReg1274_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1263_out;
SharedReg1307_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1307_out;
SharedReg332_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg332_out;
SharedReg965_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg965_out;
SharedReg1043_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1043_out;
SharedReg1133_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1133_out;
   MUX_Product310_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg103_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1293_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg965_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1043_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1133_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1039_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1094_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay102No3_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1305_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1274_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1263_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1307_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg332_out_to_MUX_Product310_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_3_impl_1_out);

   Delay1No67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_3_impl_1_out,
                 Y => Delay1No67_out);

Delay1No68_out_to_Product310_4_impl_parent_implementedSystem_port_0_cast <= Delay1No68_out;
Delay1No69_out_to_Product310_4_impl_parent_implementedSystem_port_1_cast <= Delay1No69_out;
   Product310_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_4_impl_out,
                 X => Delay1No68_out_to_Product310_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No69_out_to_Product310_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1266_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1266_out;
SharedReg666_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg666_out;
SharedReg519_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg519_out;
SharedReg614_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg614_out;
SharedReg816_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg816_out;
SharedReg520_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg520_out;
Delay87No10_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_7_cast <= Delay87No10_out;
SharedReg1305_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1305_out;
SharedReg1274_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1263_out;
SharedReg572_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg572_out;
SharedReg661_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg661_out;
SharedReg1256_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1256_out;
   MUX_Product310_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1266_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg666_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg572_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg661_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1256_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg519_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg614_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg816_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg520_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay87No10_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1305_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1274_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1263_out_to_MUX_Product310_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_4_impl_0_out);

   Delay1No68_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_4_impl_0_out,
                 Y => Delay1No68_out);

SharedReg1266_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1266_out;
SharedReg342_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg342_out;
SharedReg113_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg113_out;
SharedReg1076_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1076_out;
SharedReg1294_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1294_out;
SharedReg1271_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1271_out;
Delay102No4_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_7_cast <= Delay102No4_out;
SharedReg1305_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1305_out;
SharedReg1274_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1263_out;
SharedReg1307_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1307_out;
SharedReg341_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg341_out;
SharedReg1115_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1115_out;
   MUX_Product310_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1266_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg342_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1307_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg341_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1115_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg113_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1076_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1294_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1271_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay102No4_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1305_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1274_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1263_out_to_MUX_Product310_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_4_impl_1_out);

   Delay1No69_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_4_impl_1_out,
                 Y => Delay1No69_out);

Delay1No70_out_to_Product310_5_impl_parent_implementedSystem_port_0_cast <= Delay1No70_out;
Delay1No71_out_to_Product310_5_impl_parent_implementedSystem_port_1_cast <= Delay1No71_out;
   Product310_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product310_5_impl_out,
                 X => Delay1No70_out_to_Product310_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No71_out_to_Product310_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1264_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1264_out;
SharedReg876_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg876_out;
SharedReg1256_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1256_out;
SharedReg1266_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1266_out;
SharedReg1267_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1267_out;
SharedReg1268_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1268_out;
SharedReg1269_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1269_out;
SharedReg877_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg877_out;
SharedReg1271_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1271_out;
SharedReg1299_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1299_out;
SharedReg718_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg718_out;
SharedReg1313_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1313_out;
SharedReg1263_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1263_out;
   MUX_Product310_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1264_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg876_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg718_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1313_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1263_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1256_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1266_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1267_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1268_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1269_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg877_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1271_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1299_out_to_MUX_Product310_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_5_impl_0_out);

   Delay1No70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_5_impl_0_out,
                 Y => Delay1No70_out);

SharedReg1264_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1264_out;
Delay94No5_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_2_cast <= Delay94No5_out;
SharedReg1104_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1104_out;
SharedReg1266_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1266_out;
SharedReg1267_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1267_out;
SharedReg1268_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1268_out;
SharedReg1269_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1269_out;
SharedReg1310_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1310_out;
SharedReg1271_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1271_out;
SharedReg1299_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1299_out;
SharedReg1053_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1053_out;
SharedReg1313_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1313_out;
SharedReg1263_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1263_out;
   MUX_Product310_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1264_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay94No5_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1053_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1313_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1263_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1104_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1266_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1267_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1268_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1269_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1310_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1271_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1299_out_to_MUX_Product310_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product310_5_impl_1_out);

   Delay1No71_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product310_5_impl_1_out,
                 Y => Delay1No71_out);

Delay1No72_out_to_Product410_0_impl_parent_implementedSystem_port_0_cast <= Delay1No72_out;
Delay1No73_out_to_Product410_0_impl_parent_implementedSystem_port_1_cast <= Delay1No73_out;
   Product410_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product410_0_impl_out,
                 X => Delay1No72_out_to_Product410_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No73_out_to_Product410_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1306_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1306_out;
SharedReg300_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg300_out;
SharedReg1287_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1287_out;
SharedReg627_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg627_out;
SharedReg1256_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1256_out;
Delay78No18_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_6_cast <= Delay78No18_out;
SharedReg678_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg678_out;
SharedReg628_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg628_out;
SharedReg176_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg176_out;
SharedReg493_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg493_out;
SharedReg69_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg69_out;
SharedReg588_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg588_out;
SharedReg130_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg130_out;
   MUX_Product410_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1306_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg300_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg69_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg588_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg130_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1287_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg627_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1256_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay78No18_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg678_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg628_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg176_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg493_out_to_MUX_Product410_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_0_impl_0_out);

   Delay1No72_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_0_impl_0_out,
                 Y => Delay1No72_out);

SharedReg1306_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1306_out;
SharedReg174_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg174_out;
SharedReg1287_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1287_out;
SharedReg1277_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1277_out;
SharedReg1141_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1141_out;
SharedReg247_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg247_out;
SharedReg1317_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1317_out;
SharedReg182_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg182_out;
SharedReg240_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg240_out;
Delay78No24_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_10_cast <= Delay78No24_out;
SharedReg303_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg303_out;
SharedReg1284_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1284_out;
SharedReg304_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg304_out;
   MUX_Product410_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1306_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg174_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg303_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1284_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg304_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1287_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1277_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1141_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg247_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1317_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg182_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg240_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay78No24_out_to_MUX_Product410_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_0_impl_1_out);

   Delay1No73_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_0_impl_1_out,
                 Y => Delay1No73_out);

Delay1No74_out_to_Product410_1_impl_parent_implementedSystem_port_0_cast <= Delay1No74_out;
Delay1No75_out_to_Product410_1_impl_parent_implementedSystem_port_1_cast <= Delay1No75_out;
   Product410_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product410_1_impl_out,
                 X => Delay1No74_out_to_Product410_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No75_out_to_Product410_1_impl_parent_implementedSystem_port_1_cast);

SharedReg1272_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1272_out;
SharedReg138_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg138_out;
SharedReg1306_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1306_out;
SharedReg499_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg499_out;
SharedReg1264_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1264_out;
SharedReg1265_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1265_out;
SharedReg1256_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1256_out;
Delay78No19_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_8_cast <= Delay78No19_out;
SharedReg736_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg736_out;
SharedReg783_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg783_out;
SharedReg187_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg187_out;
SharedReg499_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg499_out;
SharedReg79_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg79_out;
   MUX_Product410_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1272_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg138_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg187_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg499_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg79_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1306_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg499_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1264_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1265_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1256_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay78No19_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg736_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg783_out_to_MUX_Product410_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_1_impl_0_out);

   Delay1No74_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_1_impl_0_out,
                 Y => Delay1No74_out);

SharedReg1272_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1272_out;
SharedReg992_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg992_out;
SharedReg1306_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1306_out;
SharedReg1275_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1275_out;
SharedReg1264_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1264_out;
SharedReg1265_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1265_out;
SharedReg1063_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1063_out;
SharedReg257_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg257_out;
SharedReg1317_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1317_out;
SharedReg193_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg193_out;
SharedReg250_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg250_out;
Delay78No25_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_12_cast <= Delay78No25_out;
SharedReg312_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg312_out;
   MUX_Product410_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1272_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg992_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg250_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay78No25_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg312_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1306_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1275_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1264_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1265_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1063_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg257_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1317_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg193_out_to_MUX_Product410_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_1_impl_1_out);

   Delay1No75_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_1_impl_1_out,
                 Y => Delay1No75_out);

Delay1No76_out_to_Product410_2_impl_parent_implementedSystem_port_0_cast <= Delay1No76_out;
Delay1No77_out_to_Product410_2_impl_parent_implementedSystem_port_1_cast <= Delay1No77_out;
   Product410_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product410_2_impl_out,
                 X => Delay1No76_out_to_Product410_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No77_out_to_Product410_2_impl_parent_implementedSystem_port_1_cast);

SharedReg463_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg463_out;
SharedReg943_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg943_out;
SharedReg1272_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1272_out;
SharedReg651_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg651_out;
SharedReg1313_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1313_out;
SharedReg1263_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1263_out;
SharedReg1264_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1264_out;
SharedReg1265_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1265_out;
SharedReg1256_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1256_out;
Delay78No20_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_10_cast <= Delay78No20_out;
SharedReg793_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg793_out;
SharedReg792_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg792_out;
SharedReg198_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg198_out;
   MUX_Product410_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg463_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg943_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg793_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg792_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg198_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1272_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg651_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1313_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1263_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1264_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1265_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1256_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay78No20_out_to_MUX_Product410_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_2_impl_0_out);

   Delay1No76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_2_impl_0_out,
                 Y => Delay1No76_out);

SharedReg145_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg145_out;
SharedReg1002_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1002_out;
SharedReg1272_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1272_out;
SharedReg1008_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1008_out;
SharedReg1313_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1313_out;
SharedReg1263_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1263_out;
SharedReg1264_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1264_out;
SharedReg1265_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1265_out;
SharedReg1022_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1022_out;
SharedReg267_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg267_out;
SharedReg1317_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1317_out;
SharedReg204_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg204_out;
SharedReg260_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg260_out;
   MUX_Product410_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg145_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1002_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1317_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg204_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg260_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1272_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1008_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1313_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1263_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1264_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1265_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1022_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg267_out_to_MUX_Product410_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_2_impl_1_out);

   Delay1No77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_2_impl_1_out,
                 Y => Delay1No77_out);

Delay1No78_out_to_Product410_3_impl_parent_implementedSystem_port_0_cast <= Delay1No78_out;
Delay1No79_out_to_Product410_3_impl_parent_implementedSystem_port_1_cast <= Delay1No79_out;
   Product410_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product410_3_impl_out,
                 X => Delay1No78_out_to_Product410_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No79_out_to_Product410_3_impl_parent_implementedSystem_port_1_cast);

SharedReg511_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg511_out;
SharedReg707_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg707_out;
SharedReg471_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg471_out;
SharedReg1127_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1127_out;
SharedReg1299_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1299_out;
SharedReg1273_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1273_out;
SharedReg1313_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1313_out;
SharedReg1263_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1263_out;
SharedReg1264_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1264_out;
SharedReg1265_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1265_out;
SharedReg1256_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1256_out;
SharedReg861_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg861_out;
SharedReg902_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg902_out;
   MUX_Product410_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg511_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg707_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1256_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg861_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg902_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg471_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1127_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1299_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1273_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1313_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1263_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1264_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1265_out_to_MUX_Product410_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_3_impl_0_out);

   Delay1No78_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_3_impl_0_out,
                 Y => Delay1No78_out);

SharedReg105_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg105_out;
SharedReg1033_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1033_out;
SharedReg153_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg153_out;
SharedReg330_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg330_out;
SharedReg1299_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1299_out;
SharedReg1273_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1273_out;
SharedReg1313_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1313_out;
SharedReg1263_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1263_out;
SharedReg1264_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1264_out;
SharedReg1265_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1265_out;
Delay9No39_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_11_cast <= Delay9No39_out;
SharedReg277_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg277_out;
SharedReg1317_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1317_out;
   MUX_Product410_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg105_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1033_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay9No39_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg277_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1317_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg153_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg330_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1299_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1273_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1313_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1263_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1264_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1265_out_to_MUX_Product410_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_3_impl_1_out);

   Delay1No79_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_3_impl_1_out,
                 Y => Delay1No79_out);

Delay1No80_out_to_Product410_4_impl_parent_implementedSystem_port_0_cast <= Delay1No80_out;
Delay1No81_out_to_Product410_4_impl_parent_implementedSystem_port_1_cast <= Delay1No81_out;
   Product410_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product410_4_impl_out,
                 X => Delay1No80_out_to_Product410_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No81_out_to_Product410_4_impl_parent_implementedSystem_port_1_cast);

SharedReg612_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg612_out;
SharedReg668_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg668_out;
SharedReg517_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg517_out;
SharedReg1293_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1293_out;
SharedReg1178_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1178_out;
SharedReg1271_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1271_out;
SharedReg1299_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1299_out;
SharedReg1273_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1273_out;
SharedReg1313_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1313_out;
SharedReg1263_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1263_out;
SharedReg1264_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1264_out;
SharedReg1265_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1265_out;
SharedReg1256_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1256_out;
   MUX_Product410_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg612_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg668_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1264_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1265_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1256_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg517_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1293_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1178_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1271_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1299_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1273_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1313_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1263_out_to_MUX_Product410_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_4_impl_0_out);

   Delay1No80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_4_impl_0_out,
                 Y => Delay1No80_out);

SharedReg1125_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1125_out;
SharedReg1075_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1075_out;
SharedReg115_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg115_out;
SharedReg1293_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1293_out;
SharedReg1310_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1310_out;
SharedReg1271_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1271_out;
SharedReg1299_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1299_out;
SharedReg1273_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1273_out;
SharedReg1313_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1313_out;
SharedReg1263_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1263_out;
SharedReg1264_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1264_out;
SharedReg1265_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1265_out;
SharedReg1119_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1119_out;
   MUX_Product410_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1125_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1075_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1264_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1265_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1119_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg115_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1293_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1310_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1271_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1299_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1273_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1313_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1263_out_to_MUX_Product410_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_4_impl_1_out);

   Delay1No81_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_4_impl_1_out,
                 Y => Delay1No81_out);

Delay1No82_out_to_Product410_5_impl_parent_implementedSystem_port_0_cast <= Delay1No82_out;
Delay1No83_out_to_Product410_5_impl_parent_implementedSystem_port_1_cast <= Delay1No83_out;
   Product410_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product410_5_impl_out,
                 X => Delay1No82_out_to_Product410_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No83_out_to_Product410_5_impl_parent_implementedSystem_port_1_cast);

SharedReg671_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg671_out;
SharedReg769_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg769_out;
SharedReg1256_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1256_out;
SharedReg526_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg526_out;
SharedReg875_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg875_out;
SharedReg626_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg626_out;
SharedReg623_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg623_out;
SharedReg1282_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1282_out;
SharedReg1104_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1104_out;
SharedReg1312_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1312_out;
SharedReg577_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg577_out;
SharedReg1274_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1263_out;
   MUX_Product410_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg671_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg769_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg577_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1274_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1263_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1256_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg526_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg875_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg626_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg623_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1282_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1104_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1312_out_to_MUX_Product410_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_5_impl_0_out);

   Delay1No82_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_5_impl_0_out,
                 Y => Delay1No82_out);

SharedReg353_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg353_out;
SharedReg1277_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1277_out;
SharedReg1109_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1109_out;
SharedReg1114_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1114_out;
SharedReg1317_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1317_out;
SharedReg64_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg64_out;
SharedReg1051_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1051_out;
SharedReg1282_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1282_out;
SharedReg1248_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1248_out;
SharedReg1312_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1312_out;
SharedReg1252_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1252_out;
SharedReg1274_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1263_out;
   MUX_Product410_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg353_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1277_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1252_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1274_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1263_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1109_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1114_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1317_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg64_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1051_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1282_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1248_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1312_out_to_MUX_Product410_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product410_5_impl_1_out);

   Delay1No83_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product410_5_impl_1_out,
                 Y => Delay1No83_out);

Delay1No84_out_to_Product510_0_impl_parent_implementedSystem_port_0_cast <= Delay1No84_out;
Delay1No85_out_to_Product510_0_impl_parent_implementedSystem_port_1_cast <= Delay1No85_out;
   Product510_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product510_0_impl_out,
                 X => Delay1No84_out_to_Product510_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No85_out_to_Product510_0_impl_parent_implementedSystem_port_1_cast);

SharedReg184_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg184_out;
SharedReg66_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg66_out;
SharedReg1264_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1264_out;
SharedReg1086_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1086_out;
SharedReg1256_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1256_out;
SharedReg776_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg776_out;
SharedReg586_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg586_out;
SharedReg1309_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1309_out;
SharedReg830_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg830_out;
SharedReg358_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg358_out;
SharedReg5_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg5_out;
Delay80No_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_12_cast <= Delay80No_out;
Delay90No_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_13_cast <= Delay90No_out;
   MUX_Product510_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg184_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg66_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg5_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay80No_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay90No_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1264_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1086_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1256_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg776_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg586_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1309_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg830_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg358_out_to_MUX_Product510_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_0_impl_0_out);

   Delay1No84_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_0_impl_0_out,
                 Y => Delay1No84_out);

Delay78No6_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_1_cast <= Delay78No6_out;
SharedReg300_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg300_out;
SharedReg1264_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1264_out;
SharedReg180_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg180_out;
SharedReg932_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg932_out;
SharedReg1316_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1316_out;
SharedReg1279_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1279_out;
SharedReg1309_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1309_out;
SharedReg1304_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1304_out;
SharedReg246_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg246_out;
SharedReg244_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg244_out;
SharedReg248_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg248_out;
SharedReg990_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg990_out;
   MUX_Product510_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay78No6_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg300_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg244_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg248_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg990_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1264_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg180_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg932_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1316_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1279_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1309_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1304_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg246_out_to_MUX_Product510_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_0_impl_1_out);

   Delay1No85_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_0_impl_1_out,
                 Y => Delay1No85_out);

Delay1No86_out_to_Product510_1_impl_parent_implementedSystem_port_0_cast <= Delay1No86_out;
Delay1No87_out_to_Product510_1_impl_parent_implementedSystem_port_1_cast <= Delay1No87_out;
   Product510_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product510_1_impl_out,
                 X => Delay1No86_out_to_Product510_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No87_out_to_Product510_1_impl_parent_implementedSystem_port_1_cast);

SharedReg640_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg640_out;
SharedReg138_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg138_out;
SharedReg195_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg195_out;
SharedReg309_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg309_out;
SharedReg501_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg501_out;
SharedReg687_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg687_out;
SharedReg1256_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1256_out;
SharedReg783_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg783_out;
SharedReg594_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg594_out;
SharedReg1309_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1309_out;
SharedReg838_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg838_out;
SharedReg411_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg411_out;
SharedReg16_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg16_out;
   MUX_Product510_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg640_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg138_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg838_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg411_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg16_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg195_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg309_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg501_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg687_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1256_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg783_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg594_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1309_out_to_MUX_Product510_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_1_impl_0_out);

   Delay1No86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_1_impl_0_out,
                 Y => Delay1No86_out);

SharedReg1284_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1284_out;
SharedReg313_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg313_out;
Delay78No7_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_3_cast <= Delay78No7_out;
SharedReg185_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg185_out;
SharedReg317_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg317_out;
Delay94No1_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_6_cast <= Delay94No1_out;
SharedReg1068_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1068_out;
SharedReg1316_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1316_out;
SharedReg1279_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1279_out;
SharedReg1309_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1309_out;
SharedReg1304_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1304_out;
SharedReg256_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg256_out;
SharedReg254_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg254_out;
   MUX_Product510_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1284_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg313_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1304_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg256_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg254_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay78No7_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg185_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg317_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay94No1_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1068_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1316_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1279_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1309_out_to_MUX_Product510_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_1_impl_1_out);

   Delay1No87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_1_impl_1_out,
                 Y => Delay1No87_out);

Delay1No88_out_to_Product510_2_impl_parent_implementedSystem_port_0_cast <= Delay1No88_out;
Delay1No89_out_to_Product510_2_impl_parent_implementedSystem_port_1_cast <= Delay1No89_out;
   Product510_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product510_2_impl_out,
                 X => Delay1No88_out_to_Product510_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No89_out_to_Product510_2_impl_parent_implementedSystem_port_1_cast);

SharedReg504_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg504_out;
SharedReg89_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg89_out;
SharedReg696_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg696_out;
SharedReg146_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg146_out;
SharedReg1274_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1263_out;
SharedReg552_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg552_out;
SharedReg694_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg694_out;
SharedReg1256_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1256_out;
SharedReg1161_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1161_out;
SharedReg646_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg646_out;
SharedReg1309_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1309_out;
SharedReg381_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg381_out;
   MUX_Product510_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg504_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg89_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg646_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1309_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg381_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg696_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg146_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1274_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1263_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg552_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg694_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1256_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1161_out_to_MUX_Product510_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_2_impl_0_out);

   Delay1No88_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_2_impl_0_out,
                 Y => Delay1No88_out);

SharedReg955_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg955_out;
SharedReg321_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg321_out;
SharedReg1284_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1284_out;
SharedReg1003_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1003_out;
SharedReg1274_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1263_out;
SharedReg326_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg326_out;
Delay94No2_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_8_cast <= Delay94No2_out;
SharedReg963_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg963_out;
SharedReg1316_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1316_out;
SharedReg1279_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1279_out;
SharedReg1309_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1309_out;
SharedReg1304_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1304_out;
   MUX_Product510_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg955_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg321_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1279_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1309_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1304_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1284_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1003_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1274_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1263_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg326_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay94No2_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg963_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1316_out_to_MUX_Product510_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_2_impl_1_out);

   Delay1No89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_2_impl_1_out,
                 Y => Delay1No89_out);

Delay1No90_out_to_Product510_3_impl_parent_implementedSystem_port_0_cast <= Delay1No90_out;
Delay1No91_out_to_Product510_3_impl_parent_implementedSystem_port_1_cast <= Delay1No91_out;
   Product510_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product510_3_impl_out,
                 X => Delay1No90_out_to_Product510_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No91_out_to_Product510_3_impl_parent_implementedSystem_port_1_cast);

SharedReg801_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg801_out;
SharedReg209_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg209_out;
SharedReg511_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg511_out;
SharedReg1127_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1127_out;
SharedReg1312_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1312_out;
SharedReg605_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg605_out;
SharedReg1274_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1263_out;
SharedReg559_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg559_out;
SharedReg759_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg759_out;
SharedReg1256_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1256_out;
SharedReg1168_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1168_out;
SharedReg704_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg704_out;
   MUX_Product510_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg801_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg209_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1256_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1168_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg704_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg511_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1127_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1312_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg605_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1274_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1263_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg559_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg759_out_to_MUX_Product510_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_3_impl_0_out);

   Delay1No90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_3_impl_0_out,
                 Y => Delay1No90_out);

SharedReg215_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg215_out;
SharedReg270_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg270_out;
Delay78No27_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_3_cast <= Delay78No27_out;
SharedReg1094_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1094_out;
SharedReg1312_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1312_out;
SharedReg1135_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1135_out;
SharedReg1274_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1263_out;
SharedReg335_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg335_out;
Delay94No3_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_10_cast <= Delay94No3_out;
SharedReg1041_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1041_out;
SharedReg1316_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1316_out;
SharedReg1279_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1279_out;
   MUX_Product510_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg215_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg270_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1041_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1316_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1279_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay78No27_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1094_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1312_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1135_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1274_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1263_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg335_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay94No3_out_to_MUX_Product510_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_3_impl_1_out);

   Delay1No91_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_3_impl_1_out,
                 Y => Delay1No91_out);

Delay1No92_out_to_Product510_4_impl_parent_implementedSystem_port_0_cast <= Delay1No92_out;
Delay1No93_out_to_Product510_4_impl_parent_implementedSystem_port_1_cast <= Delay1No93_out;
   Product510_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product510_4_impl_out,
                 X => Delay1No92_out_to_Product510_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No93_out_to_Product510_4_impl_parent_implementedSystem_port_1_cast);

SharedReg870_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg870_out;
SharedReg909_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg909_out;
SharedReg810_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg810_out;
SharedReg717_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg717_out;
SharedReg1282_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1282_out;
SharedReg1115_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1115_out;
SharedReg1312_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1312_out;
SharedReg661_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg661_out;
SharedReg1274_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1263_out;
SharedReg711_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg711_out;
SharedReg766_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg766_out;
SharedReg1256_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1256_out;
   MUX_Product510_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg870_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg909_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg711_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg766_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1256_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg810_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg717_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1282_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1115_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1312_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg661_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1274_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1263_out_to_MUX_Product510_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_4_impl_0_out);

   Delay1No92_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_4_impl_0_out,
                 Y => Delay1No92_out);

SharedReg287_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg287_out;
SharedReg1317_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1317_out;
SharedReg226_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg226_out;
SharedReg1120_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1120_out;
SharedReg1282_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1282_out;
SharedReg968_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg968_out;
SharedReg1312_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1312_out;
SharedReg1078_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1078_out;
SharedReg1274_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1274_out;
SharedReg1263_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1263_out;
SharedReg344_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg344_out;
Delay94No4_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_12_cast <= Delay94No4_out;
SharedReg1079_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1079_out;
   MUX_Product510_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg287_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1317_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg344_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay94No4_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1079_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg226_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1120_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1282_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg968_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1312_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1078_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1274_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1263_out_to_MUX_Product510_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_4_impl_1_out);

   Delay1No93_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_4_impl_1_out,
                 Y => Delay1No93_out);

Delay1No94_out_to_Product510_5_impl_parent_implementedSystem_port_0_cast <= Delay1No94_out;
Delay1No95_out_to_Product510_5_impl_parent_implementedSystem_port_1_cast <= Delay1No95_out;
   Product510_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product510_5_impl_out,
                 X => Delay1No94_out_to_Product510_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No95_out_to_Product510_5_impl_parent_implementedSystem_port_1_cast);

SharedReg718_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg718_out;
SharedReg1049_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1049_out;
SharedReg1256_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1256_out;
SharedReg826_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg826_out;
SharedReg621_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg621_out;
SharedReg490_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg490_out;
SharedReg1293_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1293_out;
SharedReg487_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg487_out;
SharedReg1044_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1044_out;
SharedReg1272_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1272_out;
SharedReg170_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg170_out;
SharedReg673_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg673_out;
SharedReg669_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg669_out;
   MUX_Product510_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg718_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1049_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg170_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg673_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg669_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1256_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg826_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg621_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg490_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1293_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg487_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1044_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1272_out_to_MUX_Product510_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_5_impl_0_out);

   Delay1No94_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_5_impl_0_out,
                 Y => Delay1No94_out);

SharedReg234_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg234_out;
SharedReg235_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg235_out;
SharedReg1056_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1056_out;
SharedReg297_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg297_out;
SharedReg351_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg351_out;
SharedReg123_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg123_out;
SharedReg1293_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1293_out;
SharedReg1112_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1112_out;
SharedReg348_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg348_out;
SharedReg1272_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1272_out;
SharedReg1249_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1249_out;
SharedReg172_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg172_out;
SharedReg1275_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1275_out;
   MUX_Product510_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg234_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg235_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1249_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg172_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1275_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1056_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg297_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg351_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg123_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1293_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1112_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg348_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1272_out_to_MUX_Product510_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product510_5_impl_1_out);

   Delay1No95_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product510_5_impl_1_out,
                 Y => Delay1No95_out);

Delay1No96_out_to_Product610_0_impl_parent_implementedSystem_port_0_cast <= Delay1No96_out;
Delay1No97_out_to_Product610_0_impl_parent_implementedSystem_port_1_cast <= Delay1No97_out;
   Product610_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_0_impl_out,
                 X => Delay1No96_out_to_Product610_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No97_out_to_Product610_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1286_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1286_out;
SharedReg1148_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1148_out;
SharedReg629_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg629_out;
SharedReg677_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg677_out;
SharedReg1256_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1256_out;
SharedReg630_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg630_out;
SharedReg731_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg731_out;
SharedReg452_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg452_out;
SharedReg68_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg68_out;
SharedReg535_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg535_out;
SharedReg1082_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1082_out;
SharedReg728_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg728_out;
SharedReg72_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg72_out;
   MUX_Product610_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1286_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1148_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1082_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg728_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg72_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg629_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg677_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1256_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg630_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg731_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg452_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg68_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg535_out_to_MUX_Product610_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product610_0_impl_0_out);

   Delay1No96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_0_impl_0_out,
                 Y => Delay1No96_out);

SharedReg1286_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1286_out;
SharedReg1275_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1275_out;
SharedReg1276_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1276_out;
SharedReg1288_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1288_out;
SharedReg929_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg929_out;
SharedReg1278_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1278_out;
SharedReg1298_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1298_out;
SharedReg2_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg2_out;
SharedReg240_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg240_out;
SharedReg1282_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1282_out;
SharedReg178_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg178_out;
SharedReg7_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg7_out;
SharedReg1145_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1145_out;
   MUX_Product610_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1286_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1275_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg178_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg7_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1145_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1276_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1288_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg929_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1278_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1298_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg2_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg240_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1282_out_to_MUX_Product610_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product610_0_impl_1_out);

   Delay1No97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_0_impl_1_out,
                 Y => Delay1No97_out);

Delay1No98_out_to_Product610_1_impl_parent_implementedSystem_port_0_cast <= Delay1No98_out;
Delay1No99_out_to_Product610_1_impl_parent_implementedSystem_port_1_cast <= Delay1No99_out;
   Product610_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_1_impl_out,
                 X => Delay1No98_out_to_Product610_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No99_out_to_Product610_1_impl_parent_implementedSystem_port_1_cast);

Delay80No1_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_1_cast <= Delay80No1_out;
Delay90No1_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_2_cast <= Delay90No1_out;
SharedReg1286_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1286_out;
SharedReg76_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg76_out;
SharedReg589_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg589_out;
SharedReg684_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg684_out;
SharedReg1256_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1256_out;
SharedReg637_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg637_out;
SharedReg743_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg743_out;
SharedReg501_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg501_out;
SharedReg78_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg78_out;
SharedReg544_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg544_out;
SharedReg933_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg933_out;
   MUX_Product610_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay80No1_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay90No1_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg78_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg544_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg933_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1286_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg76_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg589_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg684_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1256_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg637_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg743_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg501_out_to_MUX_Product610_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product610_1_impl_0_out);

   Delay1No98_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_1_impl_0_out,
                 Y => Delay1No98_out);

SharedReg258_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg258_out;
SharedReg1001_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1001_out;
SharedReg1286_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1286_out;
SharedReg309_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg309_out;
SharedReg190_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg190_out;
SharedReg1277_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1277_out;
SharedReg985_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg985_out;
SharedReg1278_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1278_out;
SharedReg1298_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1298_out;
SharedReg13_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg13_out;
SharedReg250_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg250_out;
SharedReg1282_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1282_out;
SharedReg189_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg189_out;
   MUX_Product610_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg258_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1001_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg250_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1282_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg189_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1286_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg309_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg190_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1277_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg985_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1278_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1298_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg13_out_to_MUX_Product610_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product610_1_impl_1_out);

   Delay1No99_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_1_impl_1_out,
                 Y => Delay1No99_out);

Delay1No100_out_to_Product610_2_impl_parent_implementedSystem_port_0_cast <= Delay1No100_out;
Delay1No101_out_to_Product610_2_impl_parent_implementedSystem_port_1_cast <= Delay1No101_out;
   Product610_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_2_impl_out,
                 X => Delay1No100_out_to_Product610_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No101_out_to_Product610_2_impl_parent_implementedSystem_port_1_cast);

SharedReg508_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg508_out;
SharedReg27_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg27_out;
Delay80No2_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_3_cast <= Delay80No2_out;
SharedReg146_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg146_out;
SharedReg697_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg697_out;
SharedReg550_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg550_out;
SharedReg597_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg597_out;
SharedReg746_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg746_out;
SharedReg1256_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1256_out;
SharedReg693_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg693_out;
SharedReg753_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg753_out;
SharedReg599_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg599_out;
SharedReg88_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg88_out;
   MUX_Product610_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg508_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg27_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg753_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg599_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg88_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay80No2_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg146_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg697_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg550_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg597_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg746_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1256_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg693_out_to_MUX_Product610_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product610_2_impl_0_out);

   Delay1No100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_2_impl_0_out,
                 Y => Delay1No100_out);

SharedReg266_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg266_out;
SharedReg264_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg264_out;
SharedReg268_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg268_out;
SharedReg322_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg322_out;
SharedReg148_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg148_out;
SharedReg1275_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1275_out;
SharedReg201_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg201_out;
SharedReg1277_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1277_out;
SharedReg998_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg998_out;
SharedReg1278_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1278_out;
SharedReg1298_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1298_out;
SharedReg24_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg24_out;
SharedReg260_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg260_out;
   MUX_Product610_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg266_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg264_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1298_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg24_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg260_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg268_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg322_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg148_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1275_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg201_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1277_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg998_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1278_out_to_MUX_Product610_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product610_2_impl_1_out);

   Delay1No101_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_2_impl_1_out,
                 Y => Delay1No101_out);

Delay1No102_out_to_Product610_3_impl_parent_implementedSystem_port_0_cast <= Delay1No102_out;
Delay1No103_out_to_Product610_3_impl_parent_implementedSystem_port_1_cast <= Delay1No103_out;
   Product610_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_3_impl_out,
                 X => Delay1No102_out_to_Product610_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No103_out_to_Product610_3_impl_parent_implementedSystem_port_1_cast);

SharedReg1309_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1309_out;
SharedReg390_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg390_out;
SharedReg514_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg514_out;
SharedReg99_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg99_out;
SharedReg1272_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1272_out;
SharedReg660_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg660_out;
SharedReg706_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg706_out;
SharedReg605_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg605_out;
SharedReg755_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg755_out;
SharedReg852_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg852_out;
SharedReg1256_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1256_out;
SharedReg758_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg758_out;
SharedReg807_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg807_out;
   MUX_Product610_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1309_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg390_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1256_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg758_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg807_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg514_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg99_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1272_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg660_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg706_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg605_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg755_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg852_out_to_MUX_Product610_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product610_3_impl_0_out);

   Delay1No102_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_3_impl_0_out,
                 Y => Delay1No102_out);

SharedReg1309_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1309_out;
SharedReg1304_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1304_out;
SharedReg276_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg276_out;
SharedReg330_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg330_out;
SharedReg1272_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1272_out;
SharedReg1099_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1099_out;
SharedReg156_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg156_out;
SharedReg1275_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1275_out;
SharedReg212_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg212_out;
SharedReg1277_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1277_out;
SharedReg961_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg961_out;
SharedReg1278_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1278_out;
SharedReg1298_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1298_out;
   MUX_Product610_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1309_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1304_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg961_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1278_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1298_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg276_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg330_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1272_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1099_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg156_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1275_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg212_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1277_out_to_MUX_Product610_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product610_3_impl_1_out);

   Delay1No103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_3_impl_1_out,
                 Y => Delay1No103_out);

Delay1No104_out_to_Product610_4_impl_parent_implementedSystem_port_0_cast <= Delay1No104_out;
Delay1No105_out_to_Product610_4_impl_parent_implementedSystem_port_1_cast <= Delay1No105_out;
   Product610_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_4_impl_out,
                 X => Delay1No104_out_to_Product610_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No105_out_to_Product610_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1175_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1175_out;
SharedReg812_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg812_out;
SharedReg1309_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1309_out;
SharedReg220_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg220_out;
SharedReg479_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg479_out;
SharedReg1070_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1070_out;
SharedReg1272_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1272_out;
Delay19No10_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_8_cast <= Delay19No10_out;
SharedReg715_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg715_out;
SharedReg709_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg709_out;
SharedReg762_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg762_out;
SharedReg862_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg862_out;
SharedReg1256_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1256_out;
   MUX_Product610_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1175_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg812_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg762_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg862_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1256_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1309_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg220_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg479_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1070_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1272_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay19No10_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg715_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg709_out_to_MUX_Product610_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product610_4_impl_0_out);

   Delay1No104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_4_impl_0_out,
                 Y => Delay1No104_out);

SharedReg1316_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1316_out;
SharedReg1279_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1279_out;
SharedReg1309_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1309_out;
SharedReg280_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg280_out;
SharedReg1123_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1123_out;
SharedReg339_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg339_out;
SharedReg1272_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1272_out;
SharedReg974_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg974_out;
SharedReg164_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg164_out;
SharedReg1275_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1275_out;
SharedReg223_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg223_out;
SharedReg1277_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1277_out;
SharedReg1036_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1036_out;
   MUX_Product610_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1316_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1279_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg223_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1277_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1036_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1309_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg280_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1123_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg339_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1272_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg974_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg164_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1275_out_to_MUX_Product610_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product610_4_impl_1_out);

   Delay1No105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_4_impl_1_out,
                 Y => Delay1No105_out);

Delay1No106_out_to_Product610_5_impl_parent_implementedSystem_port_0_cast <= Delay1No106_out;
Delay1No107_out_to_Product610_5_impl_parent_implementedSystem_port_1_cast <= Delay1No107_out;
   Product610_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product610_5_impl_out,
                 X => Delay1No106_out_to_Product610_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No107_out_to_Product610_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1287_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1287_out;
SharedReg873_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg873_out;
SharedReg1256_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1256_out;
SharedReg914_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg914_out;
SharedReg624_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg624_out;
SharedReg442_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg442_out;
SharedReg674_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg674_out;
SharedReg524_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg524_out;
SharedReg1044_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1044_out;
SharedReg1272_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1272_out;
SharedReg170_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg170_out;
SharedReg1306_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1306_out;
SharedReg345_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg345_out;
   MUX_Product610_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1287_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg873_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg170_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1306_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg345_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1256_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg914_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg624_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg442_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg674_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg524_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1044_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1272_out_to_MUX_Product610_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product610_5_impl_0_out);

   Delay1No106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_5_impl_0_out,
                 Y => Delay1No106_out);

SharedReg1287_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1287_out;
SharedReg1288_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1288_out;
SharedReg1015_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1015_out;
SharedReg1316_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1316_out;
SharedReg1050_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1050_out;
SharedReg125_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg125_out;
SharedReg1110_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1110_out;
SharedReg169_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg169_out;
SharedReg1248_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1248_out;
SharedReg1272_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1272_out;
SharedReg349_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg349_out;
SharedReg1306_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1306_out;
SharedReg229_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg229_out;
   MUX_Product610_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1287_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1288_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg349_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1306_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg229_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1015_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1316_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1050_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg125_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1110_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg169_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1248_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1272_out_to_MUX_Product610_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product610_5_impl_1_out);

   Delay1No107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product610_5_impl_1_out,
                 Y => Delay1No107_out);

Delay1No108_out_to_Product710_0_impl_parent_implementedSystem_port_0_cast <= Delay1No108_out;
Delay1No109_out_to_Product710_0_impl_parent_implementedSystem_port_1_cast <= Delay1No109_out;
   Product710_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product710_0_impl_out,
                 X => Delay1No108_out_to_Product710_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No109_out_to_Product710_0_impl_parent_implementedSystem_port_1_cast);

SharedReg74_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg74_out;
SharedReg1149_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1149_out;
SharedReg1085_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1085_out;
SharedReg1148_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1148_out;
SharedReg1256_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1256_out;
SharedReg1090_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1090_out;
SharedReg777_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg777_out;
SharedReg678_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg678_out;
SharedReg1088_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1088_out;
SharedReg3_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg3_out;
SharedReg729_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg729_out;
SharedReg778_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg778_out;
SharedReg986_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg986_out;
   MUX_Product710_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg74_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1149_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg729_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg778_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg986_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1085_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1148_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1256_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1090_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg777_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg678_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1088_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg3_out_to_MUX_Product710_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product710_0_impl_0_out);

   Delay1No108_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_0_impl_0_out,
                 Y => Delay1No108_out);

SharedReg249_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg249_out;
SharedReg1275_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1275_out;
SharedReg979_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg979_out;
SharedReg1277_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1277_out;
SharedReg926_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg926_out;
SharedReg1146_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1146_out;
SharedReg1296_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1296_out;
SharedReg1309_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1309_out;
SharedReg1142_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1142_out;
SharedReg129_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg129_out;
SharedReg1283_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1283_out;
SharedReg1284_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1284_out;
SharedReg133_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg133_out;
   MUX_Product710_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg249_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1275_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1283_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1284_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg133_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg979_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1277_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg926_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1146_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1296_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1309_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1142_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg129_out_to_MUX_Product710_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product710_0_impl_1_out);

   Delay1No109_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_0_impl_1_out,
                 Y => Delay1No109_out);

Delay1No110_out_to_Product710_1_impl_parent_implementedSystem_port_0_cast <= Delay1No110_out;
Delay1No111_out_to_Product710_1_impl_parent_implementedSystem_port_1_cast <= Delay1No111_out;
   Product710_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product710_1_impl_out,
                 X => Delay1No110_out_to_Product710_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No111_out_to_Product710_1_impl_parent_implementedSystem_port_1_cast);

SharedReg739_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg739_out;
SharedReg82_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg82_out;
SharedReg84_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg84_out;
SharedReg1153_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1153_out;
SharedReg1287_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1287_out;
SharedReg937_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg937_out;
SharedReg1256_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1256_out;
SharedReg942_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg942_out;
SharedReg837_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg837_out;
SharedReg686_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg686_out;
SharedReg939_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg939_out;
SharedReg14_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg14_out;
SharedReg740_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg740_out;
   MUX_Product710_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg739_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg82_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg939_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg14_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg740_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg84_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1153_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1287_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg937_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1256_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg942_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg837_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg686_out_to_MUX_Product710_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product710_1_impl_0_out);

   Delay1No110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_1_impl_0_out,
                 Y => Delay1No110_out);

SharedReg18_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg18_out;
SharedReg1067_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1067_out;
SharedReg259_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg259_out;
SharedReg1275_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1275_out;
SharedReg1287_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1287_out;
SharedReg191_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg191_out;
SharedReg945_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg945_out;
SharedReg1069_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1069_out;
SharedReg1296_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1296_out;
SharedReg1309_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1309_out;
SharedReg1064_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1064_out;
SharedReg137_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg137_out;
SharedReg1283_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1283_out;
   MUX_Product710_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg18_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1067_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1064_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg137_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1283_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg259_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1275_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1287_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg191_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg945_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1069_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1296_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1309_out_to_MUX_Product710_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product710_1_impl_1_out);

   Delay1No111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_1_impl_1_out,
                 Y => Delay1No111_out);

Delay1No112_out_to_Product710_2_impl_parent_implementedSystem_port_0_cast <= Delay1No112_out;
Delay1No113_out_to_Product710_2_impl_parent_implementedSystem_port_1_cast <= Delay1No113_out;
   Product710_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product710_2_impl_out,
                 X => Delay1No112_out_to_Product710_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No113_out_to_Product710_2_impl_parent_implementedSystem_port_1_cast);

SharedReg604_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg604_out;
SharedReg943_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg943_out;
SharedReg900_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg900_out;
Delay90No2_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_4_cast <= Delay90No2_out;
SharedReg1306_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1306_out;
SharedReg318_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg318_out;
SharedReg1287_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1287_out;
SharedReg947_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg947_out;
SharedReg1256_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1256_out;
SharedReg954_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg954_out;
SharedReg896_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg896_out;
SharedReg845_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg845_out;
SharedReg949_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg949_out;
   MUX_Product710_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg604_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg943_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg896_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg845_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg949_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg900_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay90No2_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1306_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg318_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1287_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg947_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1256_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg954_out_to_MUX_Product710_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product710_2_impl_0_out);

   Delay1No112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_2_impl_0_out,
                 Y => Delay1No112_out);

SharedReg1282_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1282_out;
SharedReg200_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg200_out;
SharedReg29_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg29_out;
SharedReg1010_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1010_out;
SharedReg1306_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1306_out;
SharedReg196_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg196_out;
SharedReg1287_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1287_out;
SharedReg202_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg202_out;
SharedReg958_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg958_out;
SharedReg1027_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1027_out;
SharedReg1296_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1296_out;
SharedReg1309_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1309_out;
SharedReg1023_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1023_out;
   MUX_Product710_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1282_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg200_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1296_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1309_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1023_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg29_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1010_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1306_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg196_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1287_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg202_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg958_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1027_out_to_MUX_Product710_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product710_2_impl_1_out);

   Delay1No113_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_2_impl_1_out,
                 Y => Delay1No113_out);

Delay1No114_out_to_Product710_3_impl_parent_implementedSystem_port_0_cast <= Delay1No114_out;
Delay1No115_out_to_Product710_3_impl_parent_implementedSystem_port_1_cast <= Delay1No115_out;
   Product710_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product710_3_impl_out,
                 X => Delay1No114_out_to_Product710_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No115_out_to_Product710_3_impl_parent_implementedSystem_port_1_cast);

SharedReg607_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg607_out;
SharedReg98_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg98_out;
SharedReg657_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg657_out;
SharedReg38_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg38_out;
SharedReg1272_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1272_out;
SharedReg154_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg154_out;
SharedReg1306_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1306_out;
SharedReg327_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg327_out;
SharedReg1287_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1287_out;
SharedReg1132_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1132_out;
SharedReg1256_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1256_out;
SharedReg1136_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1136_out;
SharedReg389_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg389_out;
   MUX_Product710_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg607_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg98_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1256_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1136_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg389_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg657_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg38_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1272_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg154_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1306_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg327_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1287_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1132_out_to_MUX_Product710_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product710_3_impl_0_out);

   Delay1No114_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_3_impl_0_out,
                 Y => Delay1No114_out);

SharedReg35_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg35_out;
SharedReg270_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg270_out;
SharedReg1282_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1282_out;
SharedReg274_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg274_out;
SharedReg1272_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1272_out;
SharedReg1095_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1095_out;
SharedReg1306_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1306_out;
SharedReg207_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg207_out;
SharedReg1287_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1287_out;
SharedReg213_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg213_out;
SharedReg1030_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1030_out;
SharedReg1043_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1043_out;
SharedReg1296_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1296_out;
   MUX_Product710_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg35_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg270_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1030_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1043_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1296_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1282_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg274_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1272_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1095_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1306_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg207_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1287_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg213_out_to_MUX_Product710_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product710_3_impl_1_out);

   Delay1No115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_3_impl_1_out,
                 Y => Delay1No115_out);

Delay1No116_out_to_Product710_4_impl_parent_implementedSystem_port_0_cast <= Delay1No116_out;
Delay1No117_out_to_Product710_4_impl_parent_implementedSystem_port_1_cast <= Delay1No117_out;
   Product710_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product710_4_impl_out,
                 X => Delay1No116_out_to_Product710_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No117_out_to_Product710_4_impl_parent_implementedSystem_port_1_cast);

SharedReg865_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg865_out;
SharedReg869_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg869_out;
SharedReg612_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg612_out;
SharedReg1195_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1195_out;
SharedReg517_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg517_out;
SharedReg1070_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1070_out;
SharedReg1272_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1272_out;
SharedReg162_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg162_out;
SharedReg1306_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1306_out;
SharedReg336_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg336_out;
SharedReg1287_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1287_out;
SharedReg1074_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1074_out;
SharedReg1256_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1256_out;
   MUX_Product710_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg865_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg869_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1287_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1074_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1256_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg612_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1195_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg517_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1070_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1272_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg162_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1306_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg336_out_to_MUX_Product710_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product710_4_impl_0_out);

   Delay1No116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_4_impl_0_out,
                 Y => Delay1No116_out);

SharedReg1278_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1278_out;
SharedReg1298_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1298_out;
SharedReg46_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg46_out;
SharedReg1304_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1304_out;
SharedReg161_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg161_out;
SharedReg968_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg968_out;
SharedReg1272_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1272_out;
SharedReg969_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg969_out;
SharedReg1306_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1306_out;
SharedReg218_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg218_out;
SharedReg1287_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1287_out;
SharedReg224_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg224_out;
SharedReg1072_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1072_out;
   MUX_Product710_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1278_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1298_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1287_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg224_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1072_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg46_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1304_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg161_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg968_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1272_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg969_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1306_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg218_out_to_MUX_Product710_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product710_4_impl_1_out);

   Delay1No117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_4_impl_1_out,
                 Y => Delay1No117_out);

Delay1No118_out_to_Product710_5_impl_parent_implementedSystem_port_0_cast <= Delay1No118_out;
Delay1No119_out_to_Product710_5_impl_parent_implementedSystem_port_1_cast <= Delay1No119_out;
   Product710_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product710_5_impl_out,
                 X => Delay1No118_out_to_Product710_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No119_out_to_Product710_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1264_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1264_out;
SharedReg1207_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1207_out;
SharedReg1256_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1256_out;
SharedReg822_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg822_out;
SharedReg821_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg821_out;
SharedReg770_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg770_out;
SharedReg231_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg231_out;
SharedReg573_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg573_out;
SharedReg119_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg119_out;
SharedReg723_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg723_out;
Delay90No5_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_11_cast <= Delay90No5_out;
SharedReg239_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg239_out;
SharedReg116_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg116_out;
   MUX_Product710_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1264_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1207_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay90No5_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg239_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg116_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1256_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg822_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg821_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg770_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg231_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg573_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg119_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg723_out_to_MUX_Product710_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product710_5_impl_0_out);

   Delay1No118_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_5_impl_0_out,
                 Y => Delay1No118_out);

SharedReg1264_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1264_out;
SharedReg1277_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1277_out;
SharedReg1117_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1117_out;
SharedReg1278_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1278_out;
SharedReg1317_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1317_out;
SharedReg237_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg237_out;
SharedReg290_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg290_out;
Delay78No29_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_8_cast <= Delay78No29_out;
SharedReg348_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg348_out;
SharedReg1284_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1284_out;
SharedReg1254_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1254_out;
Delay78No11_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_12_cast <= Delay78No11_out;
SharedReg345_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg345_out;
   MUX_Product710_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1264_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1277_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1254_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay78No11_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg345_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1117_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1278_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1317_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg237_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg290_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay78No29_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg348_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1284_out_to_MUX_Product710_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product710_5_impl_1_out);

   Delay1No119_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product710_5_impl_1_out,
                 Y => Delay1No119_out);

Delay1No120_out_to_Product810_0_impl_parent_implementedSystem_port_0_cast <= Delay1No120_out;
Delay1No121_out_to_Product810_0_impl_parent_implementedSystem_port_1_cast <= Delay1No121_out;
   Product810_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_0_impl_out,
                 X => Delay1No120_out_to_Product810_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No121_out_to_Product810_0_impl_parent_implementedSystem_port_1_cast);

SharedReg8_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg8_out;
SharedReg_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg301_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg301_out;
SharedReg781_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg781_out;
SharedReg1256_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1256_out;
SharedReg627_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg627_out;
SharedReg832_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg832_out;
SharedReg831_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg831_out;
SharedReg1088_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1088_out;
SharedReg243_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg243_out;
SharedReg778_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg778_out;
SharedReg70_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg70_out;
SharedReg1150_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1150_out;
   MUX_Product810_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg8_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg778_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg70_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1150_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg301_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg781_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1256_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg627_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg832_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg831_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1088_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg243_out_to_MUX_Product810_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product810_0_impl_0_out);

   Delay1No120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_0_impl_0_out,
                 Y => Delay1No120_out);

SharedReg245_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg245_out;
SharedReg126_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg126_out;
SharedReg127_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg127_out;
SharedReg1301_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1301_out;
SharedReg1084_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1084_out;
SharedReg1266_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1266_out;
SharedReg1291_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1291_out;
SharedReg1280_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1280_out;
SharedReg307_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg307_out;
SharedReg1143_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1143_out;
SharedReg1283_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1283_out;
SharedReg1138_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1138_out;
SharedReg1285_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1285_out;
   MUX_Product810_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg245_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg126_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1283_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1138_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1285_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg127_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1301_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1084_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1266_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1291_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1280_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg307_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1143_out_to_MUX_Product810_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product810_0_impl_1_out);

   Delay1No121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_0_impl_1_out,
                 Y => Delay1No121_out);

Delay1No122_out_to_Product810_1_impl_parent_implementedSystem_port_0_cast <= Delay1No122_out;
Delay1No123_out_to_Product810_1_impl_parent_implementedSystem_port_1_cast <= Delay1No123_out;
   Product810_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_1_impl_out,
                 X => Delay1No122_out_to_Product810_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No123_out_to_Product810_1_impl_parent_implementedSystem_port_1_cast);

SharedReg890_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg890_out;
SharedReg999_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg999_out;
SharedReg19_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg19_out;
SharedReg1154_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1154_out;
SharedReg1264_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1264_out;
SharedReg685_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg685_out;
SharedReg1256_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1256_out;
SharedReg684_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg684_out;
SharedReg839_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg839_out;
SharedReg891_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg891_out;
SharedReg939_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg939_out;
SharedReg253_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg253_out;
SharedReg1157_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1157_out;
   MUX_Product810_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg890_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg999_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg939_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg253_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1157_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg19_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1154_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1264_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg685_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1256_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg684_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg839_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg891_out_to_MUX_Product810_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product810_1_impl_0_out);

   Delay1No122_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_1_impl_0_out,
                 Y => Delay1No122_out);

SharedReg1284_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1284_out;
SharedReg141_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg141_out;
SharedReg255_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg255_out;
SharedReg1275_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1275_out;
SharedReg1264_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1264_out;
SharedReg1288_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1288_out;
SharedReg1019_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1019_out;
SharedReg1266_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1266_out;
SharedReg1291_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1291_out;
SharedReg1280_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1280_out;
SharedReg316_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg316_out;
SharedReg1065_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1065_out;
SharedReg1283_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1283_out;
   MUX_Product810_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1284_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg141_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg316_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1065_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1283_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg255_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1275_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1264_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1288_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1019_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1266_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1291_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1280_out_to_MUX_Product810_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product810_1_impl_1_out);

   Delay1No123_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_1_impl_1_out,
                 Y => Delay1No123_out);

Delay1No124_out_to_Product810_2_impl_parent_implementedSystem_port_0_cast <= Delay1No124_out;
Delay1No125_out_to_Product810_2_impl_parent_implementedSystem_port_1_cast <= Delay1No125_out;
   Product810_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_2_impl_out,
                 X => Delay1No124_out_to_Product810_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No125_out_to_Product810_2_impl_parent_implementedSystem_port_1_cast);

SharedReg25_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg25_out;
SharedReg796_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg796_out;
SharedReg897_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg897_out;
SharedReg92_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg92_out;
SharedReg206_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg206_out;
SharedReg86_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg86_out;
SharedReg1264_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1264_out;
SharedReg748_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg748_out;
SharedReg1256_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1256_out;
SharedReg791_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg791_out;
SharedReg899_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg899_out;
SharedReg898_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg898_out;
SharedReg949_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg949_out;
   MUX_Product810_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg25_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg796_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg899_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg898_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg949_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg897_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg92_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg206_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg86_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1264_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg748_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1256_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg791_out_to_MUX_Product810_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product810_2_impl_0_out);

   Delay1No124_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_2_impl_0_out,
                 Y => Delay1No124_out);

SharedReg145_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg145_out;
SharedReg1283_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1283_out;
SharedReg1284_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1284_out;
SharedReg1026_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1026_out;
Delay78No8_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_5_cast <= Delay78No8_out;
SharedReg318_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg318_out;
SharedReg1264_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1264_out;
SharedReg1288_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1288_out;
SharedReg1092_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1092_out;
SharedReg1266_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1266_out;
SharedReg1291_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1291_out;
SharedReg1280_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1280_out;
SharedReg325_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg325_out;
   MUX_Product810_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg145_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1283_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1291_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1280_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg325_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1284_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1026_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay78No8_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg318_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1264_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1288_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1092_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1266_out_to_MUX_Product810_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product810_2_impl_1_out);

   Delay1No125_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_2_impl_1_out,
                 Y => Delay1No125_out);

Delay1No126_out_to_Product810_3_impl_parent_implementedSystem_port_0_cast <= Delay1No126_out;
Delay1No127_out_to_Product810_3_impl_parent_implementedSystem_port_1_cast <= Delay1No127_out;
   Product810_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_3_impl_out,
                 X => Delay1No126_out_to_Product810_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No127_out_to_Product810_3_impl_parent_implementedSystem_port_1_cast);

SharedReg854_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg854_out;
SharedReg1134_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1134_out;
SharedReg36_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg36_out;
SharedReg1127_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1127_out;
SharedReg804_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg804_out;
SharedReg154_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg154_out;
SharedReg217_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg217_out;
SharedReg96_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg96_out;
SharedReg1264_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1264_out;
SharedReg802_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg802_out;
SharedReg1256_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1256_out;
SharedReg800_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg800_out;
SharedReg904_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg904_out;
   MUX_Product810_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg854_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1134_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1256_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg800_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg904_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg36_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1127_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg804_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg154_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg217_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg96_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1264_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg802_out_to_MUX_Product810_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product810_3_impl_0_out);

   Delay1No126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_3_impl_0_out,
                 Y => Delay1No126_out);

SharedReg1309_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1309_out;
SharedReg1033_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1033_out;
SharedReg153_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg153_out;
SharedReg211_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg211_out;
SharedReg1284_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1284_out;
SharedReg331_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg331_out;
Delay78No9_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_7_cast <= Delay78No9_out;
SharedReg327_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg327_out;
SharedReg1264_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1264_out;
SharedReg1288_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1288_out;
SharedReg1095_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1095_out;
SharedReg1266_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1266_out;
SharedReg1291_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1291_out;
   MUX_Product810_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1309_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1033_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1095_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1266_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1291_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg153_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg211_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1284_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg331_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay78No9_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg327_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1264_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1288_out_to_MUX_Product810_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product810_3_impl_1_out);

   Delay1No127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_3_impl_1_out,
                 Y => Delay1No127_out);

Delay1No128_out_to_Product810_4_impl_parent_implementedSystem_port_0_cast <= Delay1No128_out;
Delay1No129_out_to_Product810_4_impl_parent_implementedSystem_port_1_cast <= Delay1No129_out;
   Product810_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_4_impl_out,
                 X => Delay1No128_out_to_Product810_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No129_out_to_Product810_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1080_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1080_out;
SharedReg1194_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1194_out;
SharedReg864_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg864_out;
SharedReg108_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg108_out;
SharedReg566_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg566_out;
SharedReg109_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg109_out;
SharedReg814_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg814_out;
SharedReg162_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg162_out;
SharedReg228_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg228_out;
SharedReg106_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg106_out;
SharedReg1264_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1264_out;
SharedReg908_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg908_out;
SharedReg1256_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1256_out;
   MUX_Product810_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1080_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1194_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1264_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg908_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1256_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg864_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg108_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg566_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg109_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg814_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg162_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg228_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg106_out_to_MUX_Product810_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product810_4_impl_0_out);

   Delay1No128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_4_impl_0_out,
                 Y => Delay1No128_out);

SharedReg1125_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1125_out;
SharedReg1296_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1296_out;
SharedReg1309_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1309_out;
SharedReg280_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg280_out;
SharedReg1081_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1081_out;
SharedReg339_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg339_out;
SharedReg1284_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1284_out;
SharedReg340_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg340_out;
Delay78No10_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_9_cast <= Delay78No10_out;
SharedReg336_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg336_out;
SharedReg1264_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1264_out;
SharedReg1288_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1288_out;
SharedReg1117_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1117_out;
   MUX_Product810_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1125_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1296_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1264_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1288_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1117_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1309_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg280_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1081_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg339_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1284_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg340_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay78No10_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg336_out_to_MUX_Product810_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product810_4_impl_1_out);

   Delay1No129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_4_impl_1_out,
                 Y => Delay1No129_out);

Delay1No130_out_to_Product810_5_impl_parent_implementedSystem_port_0_cast <= Delay1No130_out;
Delay1No131_out_to_Product810_5_impl_parent_implementedSystem_port_1_cast <= Delay1No131_out;
   Product810_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product810_5_impl_out,
                 X => Delay1No130_out_to_Product810_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No131_out_to_Product810_5_impl_parent_implementedSystem_port_1_cast);

SharedReg821_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg821_out;
SharedReg1190_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1190_out;
SharedReg1256_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1256_out;
SharedReg1058_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1058_out;
SharedReg773_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg773_out;
SharedReg1309_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1309_out;
SharedReg1186_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1186_out;
SharedReg491_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg491_out;
SharedReg60_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg60_out;
Delay80No5_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_10_cast <= Delay80No5_out;
SharedReg122_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg122_out;
SharedReg1286_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1286_out;
SharedReg1257_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1257_out;
   MUX_Product810_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg821_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1190_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg122_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1286_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1257_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1256_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1058_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg773_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1309_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1186_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg491_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg60_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay80No5_out_to_MUX_Product810_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product810_5_impl_0_out);

   Delay1No130_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_5_impl_0_out,
                 Y => Delay1No130_out);

SharedReg1276_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1276_out;
SharedReg1301_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1301_out;
SharedReg969_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg969_out;
SharedReg1114_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1114_out;
SharedReg1279_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1279_out;
SharedReg1309_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1309_out;
SharedReg1304_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1304_out;
SharedReg296_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg296_out;
SharedReg294_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg294_out;
SharedReg298_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg298_out;
SharedReg1113_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1113_out;
SharedReg1286_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1286_out;
SharedReg1275_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1275_out;
   MUX_Product810_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1276_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1301_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1113_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1286_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1275_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg969_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1114_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1279_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1309_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1304_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg296_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg294_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg298_out_to_MUX_Product810_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product810_5_impl_1_out);

   Delay1No131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product810_5_impl_1_out,
                 Y => Delay1No131_out);

Delay1No132_out_to_Product910_0_impl_parent_implementedSystem_port_0_cast <= Delay1No132_out;
Delay1No133_out_to_Product910_0_impl_parent_implementedSystem_port_1_cast <= Delay1No133_out;
   Product910_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product910_0_impl_out,
                 X => Delay1No132_out_to_Product910_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No133_out_to_Product910_0_impl_parent_implementedSystem_port_1_cast);

SharedReg882_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg882_out;
Delay1No332_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_2_cast <= Delay1No332_out;
SharedReg833_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg833_out;
SharedReg834_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg834_out;
SharedReg1256_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1256_out;
SharedReg1149_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1149_out;
SharedReg365_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg365_out;
SharedReg730_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg730_out;
SharedReg68_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg68_out;
SharedReg1150_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1150_out;
Delay64No_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_11_cast <= Delay64No_out;
SharedReg827_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg827_out;
SharedReg414_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg414_out;
   MUX_Product910_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg882_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No332_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay64No_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg827_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg414_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg833_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg834_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1256_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1149_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg365_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg730_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg68_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1150_out_to_MUX_Product910_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product910_0_impl_0_out);

   Delay1No132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_0_impl_0_out,
                 Y => Delay1No132_out);

SharedReg1295_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1295_out;
SharedReg1263_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1263_out;
SharedReg1276_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1276_out;
SharedReg1297_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1297_out;
SharedReg925_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg925_out;
SharedReg1290_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1290_out;
SharedReg1279_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1279_out;
SharedReg1303_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1303_out;
SharedReg128_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg128_out;
SharedReg1294_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1294_out;
SharedReg1311_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1311_out;
SharedReg1284_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1284_out;
SharedReg1305_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1305_out;
   MUX_Product910_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1295_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1263_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1311_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1284_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1305_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1276_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1297_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg925_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1290_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1279_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1303_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg128_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1294_out_to_MUX_Product910_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product910_0_impl_1_out);

   Delay1No133_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_0_impl_1_out,
                 Y => Delay1No133_out);

Delay1No134_out_to_Product910_1_impl_parent_implementedSystem_port_0_cast <= Delay1No134_out;
Delay1No135_out_to_Product910_1_impl_parent_implementedSystem_port_1_cast <= Delay1No135_out;
   Product910_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product910_1_impl_out,
                 X => Delay1No134_out_to_Product910_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No135_out_to_Product910_1_impl_parent_implementedSystem_port_1_cast);

SharedReg80_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg80_out;
SharedReg1155_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1155_out;
SharedReg890_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg890_out;
SharedReg11_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg11_out;
SharedReg636_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg636_out;
SharedReg371_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg371_out;
SharedReg1256_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1256_out;
SharedReg1154_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1154_out;
SharedReg373_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg373_out;
SharedReg741_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg741_out;
SharedReg78_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg78_out;
SharedReg420_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg420_out;
SharedReg842_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg842_out;
   MUX_Product910_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg80_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1155_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg78_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg420_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg842_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg890_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg11_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg636_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg371_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1256_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1154_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg373_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg741_out_to_MUX_Product910_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product910_1_impl_0_out);

   Delay1No134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_1_impl_0_out,
                 Y => Delay1No134_out);

SharedReg1060_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1060_out;
SharedReg1285_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1285_out;
SharedReg1295_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1295_out;
SharedReg134_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg134_out;
SharedReg1276_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1276_out;
SharedReg1277_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1277_out;
SharedReg1060_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1060_out;
SharedReg1290_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1290_out;
SharedReg1279_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1279_out;
SharedReg1303_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1303_out;
SharedReg136_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg136_out;
SharedReg1294_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1294_out;
SharedReg1311_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1311_out;
   MUX_Product910_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1060_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1285_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg136_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1294_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1311_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1295_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg134_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1276_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1277_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1060_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1290_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1279_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1303_out_to_MUX_Product910_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product910_1_impl_1_out);

   Delay1No135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_1_impl_1_out,
                 Y => Delay1No135_out);

Delay1No136_out_to_Product910_2_impl_parent_implementedSystem_port_0_cast <= Delay1No136_out;
Delay1No137_out_to_Product910_2_impl_parent_implementedSystem_port_1_cast <= Delay1No137_out;
   Product910_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product910_2_impl_out,
                 X => Delay1No136_out_to_Product910_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No137_out_to_Product910_2_impl_parent_implementedSystem_port_1_cast);

SharedReg263_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg263_out;
SharedReg1164_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1164_out;
SharedReg90_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg90_out;
SharedReg1009_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1009_out;
SharedReg1286_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1286_out;
SharedReg379_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg379_out;
SharedReg645_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg645_out;
SharedReg425_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg425_out;
SharedReg1256_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1256_out;
SharedReg472_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg472_out;
SharedReg512_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg512_out;
SharedReg752_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg752_out;
SharedReg88_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg88_out;
   MUX_Product910_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg263_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1164_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg512_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg752_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg88_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg90_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1009_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1286_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg379_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg645_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg425_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1256_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg472_out_to_MUX_Product910_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product910_2_impl_0_out);

   Delay1No136_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_2_impl_0_out,
                 Y => Delay1No136_out);

SharedReg1024_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1024_out;
SharedReg1283_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1283_out;
SharedReg1018_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1018_out;
SharedReg149_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg149_out;
SharedReg1286_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1286_out;
SharedReg1275_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1275_out;
SharedReg1276_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1276_out;
SharedReg1277_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1277_out;
SharedReg1018_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1018_out;
SharedReg1290_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1290_out;
SharedReg1279_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1279_out;
SharedReg1303_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1303_out;
SharedReg144_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg144_out;
   MUX_Product910_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1024_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1283_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1279_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1303_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg144_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1018_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg149_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1286_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1275_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1276_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1277_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1018_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1290_out_to_MUX_Product910_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product910_2_impl_1_out);

   Delay1No137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_2_impl_1_out,
                 Y => Delay1No137_out);

Delay1No138_out_to_Product910_3_impl_parent_implementedSystem_port_0_cast <= Delay1No138_out;
Delay1No139_out_to_Product910_3_impl_parent_implementedSystem_port_1_cast <= Delay1No139_out;
   Product910_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product910_3_impl_out,
                 X => Delay1No138_out_to_Product910_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No139_out_to_Product910_3_impl_parent_implementedSystem_port_1_cast);

SharedReg438_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg438_out;
SharedReg1134_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1134_out;
SharedReg273_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg273_out;
SharedReg858_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg858_out;
Delay80No3_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_5_cast <= Delay80No3_out;
Delay90No3_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_6_cast <= Delay90No3_out;
SharedReg1286_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1286_out;
SharedReg433_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg433_out;
SharedReg703_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg703_out;
SharedReg517_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg517_out;
SharedReg1256_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1256_out;
SharedReg480_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg480_out;
SharedReg518_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg518_out;
   MUX_Product910_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg438_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1134_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1256_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg480_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg518_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg273_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg858_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay80No3_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay90No3_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1286_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg433_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg703_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg517_out_to_MUX_Product910_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product910_3_impl_0_out);

   Delay1No138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_3_impl_0_out,
                 Y => Delay1No138_out);

SharedReg1280_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1280_out;
SharedReg334_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg334_out;
SharedReg1034_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1034_out;
SharedReg1283_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1283_out;
SharedReg278_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg278_out;
SharedReg1103_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1103_out;
SharedReg1286_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1286_out;
SharedReg1275_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1275_out;
SharedReg1276_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1276_out;
SharedReg1277_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1277_out;
SharedReg1128_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1128_out;
SharedReg1290_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1290_out;
SharedReg1279_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1279_out;
   MUX_Product910_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1280_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg334_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1128_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1290_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1279_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1034_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1283_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg278_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1103_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1286_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1275_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1276_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1277_out_to_MUX_Product910_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product910_3_impl_1_out);

   Delay1No139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_3_impl_1_out,
                 Y => Delay1No139_out);

Delay1No140_out_to_Product910_4_impl_parent_implementedSystem_port_0_cast <= Delay1No140_out;
Delay1No141_out_to_Product910_4_impl_parent_implementedSystem_port_1_cast <= Delay1No141_out;
   Product910_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product910_4_impl_out,
                 X => Delay1No140_out_to_Product910_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No141_out_to_Product910_4_impl_parent_implementedSystem_port_1_cast);

SharedReg809_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg809_out;
SharedReg399_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg399_out;
SharedReg398_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg398_out;
SharedReg1076_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1076_out;
SharedReg520_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg520_out;
SharedReg49_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg49_out;
Delay80No4_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_7_cast <= Delay80No4_out;
Delay90No4_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_8_cast <= Delay90No4_out;
SharedReg1286_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1286_out;
SharedReg487_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg487_out;
SharedReg764_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg764_out;
SharedReg487_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg487_out;
SharedReg1256_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1256_out;
   MUX_Product910_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg809_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg399_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg764_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg487_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1256_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg398_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1076_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg520_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg49_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay80No4_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay90No4_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1286_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg487_out_to_MUX_Product910_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product910_4_impl_0_out);

   Delay1No140_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_4_impl_0_out,
                 Y => Delay1No140_out);

SharedReg1266_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1266_out;
SharedReg1291_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1291_out;
SharedReg1280_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1280_out;
SharedReg1120_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1120_out;
SharedReg286_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg286_out;
SharedReg284_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg284_out;
SharedReg288_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg288_out;
SharedReg976_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg976_out;
SharedReg1286_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1286_out;
SharedReg1275_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1275_out;
SharedReg1276_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1276_out;
SharedReg1277_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1277_out;
SharedReg966_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg966_out;
   MUX_Product910_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1266_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1291_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1276_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1277_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg966_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1280_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1120_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg286_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg284_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg288_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg976_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1286_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1275_out_to_MUX_Product910_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product910_4_impl_1_out);

   Delay1No141_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_4_impl_1_out,
                 Y => Delay1No141_out);

Delay1No142_out_to_Product910_5_impl_parent_implementedSystem_port_0_cast <= Delay1No142_out;
Delay1No143_out_to_Product910_5_impl_parent_implementedSystem_port_1_cast <= Delay1No143_out;
   Product910_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product910_5_impl_out,
                 X => Delay1No142_out_to_Product910_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No143_out_to_Product910_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1048_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1048_out;
SharedReg1206_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1206_out;
SharedReg1256_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1256_out;
SharedReg769_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg769_out;
SharedReg921_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg921_out;
SharedReg575_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg575_out;
SharedReg118_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg118_out;
SharedReg723_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg723_out;
SharedReg1044_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1044_out;
SharedReg878_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg878_out;
SharedReg1253_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1253_out;
SharedReg124_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg124_out;
SharedReg1258_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg1258_out;
   MUX_Product910_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1048_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1206_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1253_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg124_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1258_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1256_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg769_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg921_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg575_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg118_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg723_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1044_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg878_out_to_MUX_Product910_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product910_5_impl_0_out);

   Delay1No142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_5_impl_0_out,
                 Y => Delay1No142_out);

SharedReg1250_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1250_out;
SharedReg1297_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1297_out;
SharedReg1012_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1012_out;
SharedReg1266_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1266_out;
SharedReg1298_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1298_out;
SharedReg57_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg57_out;
SharedReg290_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg290_out;
SharedReg1282_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1282_out;
SharedReg233_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg233_out;
SharedReg62_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg62_out;
SharedReg173_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg173_out;
SharedReg299_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg299_out;
SharedReg1275_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1275_out;
   MUX_Product910_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1250_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1297_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg173_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg299_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1275_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1012_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1266_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1298_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg57_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg290_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1282_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg233_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg62_out_to_MUX_Product910_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product910_5_impl_1_out);

   Delay1No143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product910_5_impl_1_out,
                 Y => Delay1No143_out);
   Inv_11_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_11_0_IEEE,
                 X => Delay1No144_out);
Inv_11_0 <= Inv_11_0_IEEE;

   Delay1No144_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg354_out,
                 Y => Delay1No144_out);
   Inv_11_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_11_1_IEEE,
                 X => Delay1No145_out);
Inv_11_1 <= Inv_11_1_IEEE;

   Delay1No145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg363_out,
                 Y => Delay1No145_out);
   Inv_11_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_11_2_IEEE,
                 X => Delay1No146_out);
Inv_11_2 <= Inv_11_2_IEEE;

   Delay1No146_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg371_out,
                 Y => Delay1No146_out);
   Inv_11_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_11_3_IEEE,
                 X => Delay1No147_out);
Inv_11_3 <= Inv_11_3_IEEE;

   Delay1No147_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg379_out,
                 Y => Delay1No147_out);
   Inv_11_4_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_11_4_IEEE,
                 X => Delay1No148_out);
Inv_11_4 <= Inv_11_4_IEEE;

   Delay1No148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg386_out,
                 Y => Delay1No148_out);
   Inv_11_5_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_11_5_IEEE,
                 X => Delay1No149_out);
Inv_11_5 <= Inv_11_5_IEEE;

   Delay1No149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg394_out,
                 Y => Delay1No149_out);
   Inv_12_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_12_0_IEEE,
                 X => Delay1No150_out);
Inv_12_0 <= Inv_12_0_IEEE;

   Delay1No150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg400_out,
                 Y => Delay1No150_out);
   Inv_12_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_12_1_IEEE,
                 X => Delay1No151_out);
Inv_12_1 <= Inv_12_1_IEEE;

   Delay1No151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg408_out,
                 Y => Delay1No151_out);
   Inv_12_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_12_2_IEEE,
                 X => Delay1No152_out);
Inv_12_2 <= Inv_12_2_IEEE;

   Delay1No152_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg418_out,
                 Y => Delay1No152_out);
   Inv_12_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_12_3_IEEE,
                 X => Delay1No153_out);
Inv_12_3 <= Inv_12_3_IEEE;

   Delay1No153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg425_out,
                 Y => Delay1No153_out);
   Inv_12_4_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_12_4_IEEE,
                 X => Delay1No154_out);
Inv_12_4 <= Inv_12_4_IEEE;

   Delay1No154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg433_out,
                 Y => Delay1No154_out);
   Inv_12_5_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_12_5_IEEE,
                 X => Delay1No155_out);
Inv_12_5 <= Inv_12_5_IEEE;

   Delay1No155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg442_out,
                 Y => Delay1No155_out);
   Inv_13_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_13_0_IEEE,
                 X => Delay1No156_out);
Inv_13_0 <= Inv_13_0_IEEE;

   Delay1No156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg531_out,
                 Y => Delay1No156_out);
   Inv_13_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_13_1_IEEE,
                 X => Delay1No157_out);
Inv_13_1 <= Inv_13_1_IEEE;

   Delay1No157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg540_out,
                 Y => Delay1No157_out);
   Inv_13_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_13_2_IEEE,
                 X => Delay1No158_out);
Inv_13_2 <= Inv_13_2_IEEE;

   Delay1No158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg550_out,
                 Y => Delay1No158_out);
   Inv_13_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_13_3_IEEE,
                 X => Delay1No159_out);
Inv_13_3 <= Inv_13_3_IEEE;

   Delay1No159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg557_out,
                 Y => Delay1No159_out);
   Inv_13_4_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_13_4_IEEE,
                 X => Delay1No160_out);
Inv_13_4 <= Inv_13_4_IEEE;

   Delay1No160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg566_out,
                 Y => Delay1No160_out);
   Inv_13_5_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_13_5_IEEE,
                 X => Delay1No161_out);
Inv_13_5 <= Inv_13_5_IEEE;

   Delay1No161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg573_out,
                 Y => Delay1No161_out);
   Inv_21_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_21_0_IEEE,
                 X => Delay1No162_out);
Inv_21_0 <= Inv_21_0_IEEE;

   Delay1No162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg581_out,
                 Y => Delay1No162_out);
   Inv_21_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_21_1_IEEE,
                 X => Delay1No163_out);
Inv_21_1 <= Inv_21_1_IEEE;

   Delay1No163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg589_out,
                 Y => Delay1No163_out);
   Inv_21_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_21_2_IEEE,
                 X => Delay1No164_out);
Inv_21_2 <= Inv_21_2_IEEE;

   Delay1No164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg597_out,
                 Y => Delay1No164_out);
   Inv_21_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_21_3_IEEE,
                 X => Delay1No165_out);
Inv_21_3 <= Inv_21_3_IEEE;

   Delay1No165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg605_out,
                 Y => Delay1No165_out);
   Inv_21_4_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_21_4_IEEE,
                 X => Delay1No166_out);
Inv_21_4 <= Inv_21_4_IEEE;

   Delay1No166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg610_out,
                 Y => Delay1No166_out);
   Inv_21_5_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_21_5_IEEE,
                 X => Delay1No167_out);
Inv_21_5 <= Inv_21_5_IEEE;

   Delay1No167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg618_out,
                 Y => Delay1No167_out);
   Inv_22_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_22_0_IEEE,
                 X => Delay1No168_out);
Inv_22_0 <= Inv_22_0_IEEE;

   Delay1No168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg627_out,
                 Y => Delay1No168_out);
   Inv_22_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_22_1_IEEE,
                 X => Delay1No169_out);
Inv_22_1 <= Inv_22_1_IEEE;

   Delay1No169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg634_out,
                 Y => Delay1No169_out);
   Inv_22_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_22_2_IEEE,
                 X => Delay1No170_out);
Inv_22_2 <= Inv_22_2_IEEE;

   Delay1No170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg642_out,
                 Y => Delay1No170_out);
   Inv_22_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_22_3_IEEE,
                 X => Delay1No171_out);
Inv_22_3 <= Inv_22_3_IEEE;

   Delay1No171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg652_out,
                 Y => Delay1No171_out);
   Inv_22_4_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_22_4_IEEE,
                 X => Delay1No172_out);
Inv_22_4 <= Inv_22_4_IEEE;

   Delay1No172_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg661_out,
                 Y => Delay1No172_out);
   Inv_22_5_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_22_5_IEEE,
                 X => Delay1No173_out);
Inv_22_5 <= Inv_22_5_IEEE;

   Delay1No173_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg669_out,
                 Y => Delay1No173_out);
   Inv_23_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_23_0_IEEE,
                 X => Delay1No174_out);
Inv_23_0 <= Inv_23_0_IEEE;

   Delay1No174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg676_out,
                 Y => Delay1No174_out);
   Inv_23_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_23_1_IEEE,
                 X => Delay1No175_out);
Inv_23_1 <= Inv_23_1_IEEE;

   Delay1No175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg684_out,
                 Y => Delay1No175_out);
   Inv_23_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_23_2_IEEE,
                 X => Delay1No176_out);
Inv_23_2 <= Inv_23_2_IEEE;

   Delay1No176_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg690_out,
                 Y => Delay1No176_out);
   Inv_23_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_23_3_IEEE,
                 X => Delay1No177_out);
Inv_23_3 <= Inv_23_3_IEEE;

   Delay1No177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg700_out,
                 Y => Delay1No177_out);
   Inv_23_4_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_23_4_IEEE,
                 X => Delay1No178_out);
Inv_23_4 <= Inv_23_4_IEEE;

   Delay1No178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg709_out,
                 Y => Delay1No178_out);
   Inv_23_5_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_23_5_IEEE,
                 X => Delay1No179_out);
Inv_23_5 <= Inv_23_5_IEEE;

   Delay1No179_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg718_out,
                 Y => Delay1No179_out);
   Inv_31_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_31_0_IEEE,
                 X => Delay1No180_out);
Inv_31_0 <= Inv_31_0_IEEE;

   Delay1No180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg726_out,
                 Y => Delay1No180_out);
   Inv_31_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_31_1_IEEE,
                 X => Delay1No181_out);
Inv_31_1 <= Inv_31_1_IEEE;

   Delay1No181_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg735_out,
                 Y => Delay1No181_out);
   Inv_31_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_31_2_IEEE,
                 X => Delay1No182_out);
Inv_31_2 <= Inv_31_2_IEEE;

   Delay1No182_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg746_out,
                 Y => Delay1No182_out);
   Inv_31_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_31_3_IEEE,
                 X => Delay1No183_out);
Inv_31_3 <= Inv_31_3_IEEE;

   Delay1No183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg755_out,
                 Y => Delay1No183_out);
   Inv_31_4_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_31_4_IEEE,
                 X => Delay1No184_out);
Inv_31_4 <= Inv_31_4_IEEE;

   Delay1No184_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg762_out,
                 Y => Delay1No184_out);
   Inv_31_5_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_31_5_IEEE,
                 X => Delay1No185_out);
Inv_31_5 <= Inv_31_5_IEEE;

   Delay1No185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg769_out,
                 Y => Delay1No185_out);
   Inv_32_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_32_0_IEEE,
                 X => Delay1No186_out);
Inv_32_0 <= Inv_32_0_IEEE;

   Delay1No186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg775_out,
                 Y => Delay1No186_out);
   Inv_32_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_32_1_IEEE,
                 X => Delay1No187_out);
Inv_32_1 <= Inv_32_1_IEEE;

   Delay1No187_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg782_out,
                 Y => Delay1No187_out);
   Inv_32_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_32_2_IEEE,
                 X => Delay1No188_out);
Inv_32_2 <= Inv_32_2_IEEE;

   Delay1No188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg791_out,
                 Y => Delay1No188_out);
   Inv_32_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_32_3_IEEE,
                 X => Delay1No189_out);
Inv_32_3 <= Inv_32_3_IEEE;

   Delay1No189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg800_out,
                 Y => Delay1No189_out);
   Inv_32_4_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_32_4_IEEE,
                 X => Delay1No190_out);
Inv_32_4 <= Inv_32_4_IEEE;

   Delay1No190_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg809_out,
                 Y => Delay1No190_out);
   Inv_32_5_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_32_5_IEEE,
                 X => Delay1No191_out);
Inv_32_5 <= Inv_32_5_IEEE;

   Delay1No191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg819_out,
                 Y => Delay1No191_out);
   Inv_33_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_33_0_IEEE,
                 X => Delay1No192_out);
Inv_33_0 <= Inv_33_0_IEEE;

   Delay1No192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg827_out,
                 Y => Delay1No192_out);
   Inv_33_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_33_1_IEEE,
                 X => Delay1No193_out);
Inv_33_1 <= Inv_33_1_IEEE;

   Delay1No193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg835_out,
                 Y => Delay1No193_out);
   Inv_33_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_33_2_IEEE,
                 X => Delay1No194_out);
Inv_33_2 <= Inv_33_2_IEEE;

   Delay1No194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg843_out,
                 Y => Delay1No194_out);
   Inv_33_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_33_3_IEEE,
                 X => Delay1No195_out);
Inv_33_3 <= Inv_33_3_IEEE;

   Delay1No195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg852_out,
                 Y => Delay1No195_out);
   Inv_33_4_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_33_4_IEEE,
                 X => Delay1No196_out);
Inv_33_4 <= Inv_33_4_IEEE;

   Delay1No196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg862_out,
                 Y => Delay1No196_out);
   Inv_33_5_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_33_5_IEEE,
                 X => Delay1No197_out);
Inv_33_5 <= Inv_33_5_IEEE;

   Delay1No197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg871_out,
                 Y => Delay1No197_out);
   Inv_41_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_41_0_IEEE,
                 X => Delay1No198_out);
Inv_41_0 <= Inv_41_0_IEEE;

   Delay1No198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg879_out,
                 Y => Delay1No198_out);
   Inv_41_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_41_1_IEEE,
                 X => Delay1No199_out);
Inv_41_1 <= Inv_41_1_IEEE;

   Delay1No199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg887_out,
                 Y => Delay1No199_out);
   Inv_41_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_41_2_IEEE,
                 X => Delay1No200_out);
Inv_41_2 <= Inv_41_2_IEEE;

   Delay1No200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg893_out,
                 Y => Delay1No200_out);
   Inv_41_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_41_3_IEEE,
                 X => Delay1No201_out);
Inv_41_3 <= Inv_41_3_IEEE;

   Delay1No201_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg901_out,
                 Y => Delay1No201_out);
   Inv_41_4_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_41_4_IEEE,
                 X => Delay1No202_out);
Inv_41_4 <= Inv_41_4_IEEE;

   Delay1No202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg907_out,
                 Y => Delay1No202_out);
   Inv_41_5_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_41_5_IEEE,
                 X => Delay1No203_out);
Inv_41_5 <= Inv_41_5_IEEE;

   Delay1No203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg913_out,
                 Y => Delay1No203_out);
   Inv_42_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_42_0_IEEE,
                 X => Delay1No204_out);
Inv_42_0 <= Inv_42_0_IEEE;

   Delay1No204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg450_out,
                 Y => Delay1No204_out);
   Inv_42_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_42_1_IEEE,
                 X => Delay1No205_out);
Inv_42_1 <= Inv_42_1_IEEE;

   Delay1No205_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg456_out,
                 Y => Delay1No205_out);
   Inv_42_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_42_2_IEEE,
                 X => Delay1No206_out);
Inv_42_2 <= Inv_42_2_IEEE;

   Delay1No206_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg463_out,
                 Y => Delay1No206_out);
   Inv_42_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_42_3_IEEE,
                 X => Delay1No207_out);
Inv_42_3 <= Inv_42_3_IEEE;

   Delay1No207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg471_out,
                 Y => Delay1No207_out);
   Inv_42_4_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_42_4_IEEE,
                 X => Delay1No208_out);
Inv_42_4 <= Inv_42_4_IEEE;

   Delay1No208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg479_out,
                 Y => Delay1No208_out);
   Inv_42_5_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_42_5_IEEE,
                 X => Delay1No209_out);
Inv_42_5 <= Inv_42_5_IEEE;

   Delay1No209_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg487_out,
                 Y => Delay1No209_out);
   Inv_43_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_43_0_IEEE,
                 X => Delay1No210_out);
Inv_43_0 <= Inv_43_0_IEEE;

   Delay1No210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg493_out,
                 Y => Delay1No210_out);
   Inv_43_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_43_1_IEEE,
                 X => Delay1No211_out);
Inv_43_1 <= Inv_43_1_IEEE;

   Delay1No211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg499_out,
                 Y => Delay1No211_out);
   Inv_43_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_43_2_IEEE,
                 X => Delay1No212_out);
Inv_43_2 <= Inv_43_2_IEEE;

   Delay1No212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg504_out,
                 Y => Delay1No212_out);
   Inv_43_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_43_3_IEEE,
                 X => Delay1No213_out);
Inv_43_3 <= Inv_43_3_IEEE;

   Delay1No213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg511_out,
                 Y => Delay1No213_out);
   Inv_43_4_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_43_4_IEEE,
                 X => Delay1No214_out);
Inv_43_4 <= Inv_43_4_IEEE;

   Delay1No214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg517_out,
                 Y => Delay1No214_out);
   Inv_43_5_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Inv_43_5_IEEE,
                 X => Delay1No215_out);
Inv_43_5 <= Inv_43_5_IEEE;

   Delay1No215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg524_out,
                 Y => Delay1No215_out);

Delay1No216_out_to_Add30_0_impl_parent_implementedSystem_port_0_cast <= Delay1No216_out;
Delay1No217_out_to_Add30_0_impl_parent_implementedSystem_port_1_cast <= Delay1No217_out;
   Add30_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_0_impl_out,
                 X => Delay1No216_out_to_Add30_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No217_out_to_Add30_0_impl_parent_implementedSystem_port_1_cast);

SharedReg633_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg633_out;
SharedReg585_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg585_out;
SharedReg400_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg400_out;
SharedReg403_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg403_out;
SharedReg356_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg356_out;
SharedReg886_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg886_out;
SharedReg582_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg582_out;
SharedReg450_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg450_out;
SharedReg363_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg363_out;
SharedReg498_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg498_out;
Delay73No6_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_11_cast <= Delay73No6_out;
Delay88No6_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_12_cast <= Delay88No6_out;
SharedReg584_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg584_out;
   MUX_Add30_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg633_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg585_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay73No6_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay88No6_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg584_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg400_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg403_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg356_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg886_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg582_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg450_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg363_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg498_out_to_MUX_Add30_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_0_impl_0_out);

   Delay1No216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_0_impl_0_out,
                 Y => Delay1No216_out);

SharedReg930_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg930_out;
SharedReg583_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg583_out;
Delay96No_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_3_cast <= Delay96No_out;
SharedReg531_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg531_out;
Delay70No_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_5_cast <= Delay70No_out;
SharedReg933_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg933_out;
SharedReg726_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg726_out;
SharedReg584_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg584_out;
SharedReg494_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg494_out;
SharedReg1217_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1217_out;
SharedReg1215_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1215_out;
SharedReg1086_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1086_out;
SharedReg1214_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1214_out;
   MUX_Add30_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg930_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg583_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1215_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1086_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1214_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay96No_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg531_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay70No_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg933_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg726_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg584_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg494_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1217_out_to_MUX_Add30_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_0_impl_1_out);

   Delay1No217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_0_impl_1_out,
                 Y => Delay1No217_out);

Delay1No218_out_to_Add30_1_impl_parent_implementedSystem_port_0_cast <= Delay1No218_out;
Delay1No219_out_to_Add30_1_impl_parent_implementedSystem_port_1_cast <= Delay1No219_out;
   Add30_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_1_impl_out,
                 X => Delay1No218_out_to_Add30_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No219_out_to_Add30_1_impl_parent_implementedSystem_port_1_cast);

SharedReg369_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg369_out;
SharedReg416_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg416_out;
SharedReg502_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg502_out;
SharedReg1155_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1155_out;
SharedReg456_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg456_out;
SharedReg459_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg459_out;
SharedReg639_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg639_out;
Delay5No1_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_8_cast <= Delay5No1_out;
SharedReg463_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg463_out;
Delay88No1_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_10_cast <= Delay88No1_out;
SharedReg422_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg422_out;
SharedReg885_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg885_out;
SharedReg532_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg532_out;
   MUX_Add30_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg369_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg416_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg422_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg885_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg532_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg502_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1155_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg456_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg459_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg639_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay5No1_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg463_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay88No1_out_to_MUX_Add30_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_1_impl_0_out);

   Delay1No218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_1_impl_0_out,
                 Y => Delay1No218_out);

SharedReg1137_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1137_out;
SharedReg933_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg933_out;
SharedReg1220_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1220_out;
SharedReg991_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg991_out;
Delay96No1_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_5_cast <= Delay96No1_out;
SharedReg589_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg589_out;
SharedReg1221_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1221_out;
SharedReg1153_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1153_out;
SharedReg1059_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1059_out;
SharedReg1219_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1219_out;
SharedReg641_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg641_out;
SharedReg1137_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1137_out;
SharedReg1215_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1215_out;
   MUX_Add30_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1137_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg933_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg641_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1137_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1215_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1220_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg991_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay96No1_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg589_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1221_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1153_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1059_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1219_out_to_MUX_Add30_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_1_impl_1_out);

   Delay1No219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_1_impl_1_out,
                 Y => Delay1No219_out);

Delay1No220_out_to_Add30_2_impl_parent_implementedSystem_port_0_cast <= Delay1No220_out;
Delay1No221_out_to_Add30_2_impl_parent_implementedSystem_port_1_cast <= Delay1No221_out;
   Add30_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_2_impl_out,
                 X => Delay1No220_out_to_Add30_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No221_out_to_Add30_2_impl_parent_implementedSystem_port_1_cast);

SharedReg738_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg738_out;
SharedReg541_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg541_out;
SharedReg466_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg466_out;
SharedReg470_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg470_out;
SharedReg754_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg754_out;
SharedReg601_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg601_out;
SharedReg463_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg463_out;
SharedReg554_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg554_out;
SharedReg648_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg648_out;
Delay5No2_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_10_cast <= Delay5No2_out;
SharedReg471_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg471_out;
SharedReg841_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg841_out;
SharedReg548_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg548_out;
   MUX_Add30_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg738_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg541_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg471_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg841_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg548_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg466_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg470_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg754_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg601_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg463_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg554_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg648_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay5No2_out_to_MUX_Add30_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_2_impl_0_out);

   Delay1No220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_2_impl_0_out,
                 Y => Delay1No220_out);

SharedReg1156_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1156_out;
SharedReg1221_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1221_out;
SharedReg1059_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1059_out;
SharedReg1002_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1002_out;
SharedReg1000_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1000_out;
SharedReg599_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg599_out;
Delay96No2_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_7_cast <= Delay96No2_out;
SharedReg642_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg642_out;
SharedReg1227_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1227_out;
SharedReg425_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg425_out;
SharedReg1002_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1002_out;
SharedReg991_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg991_out;
SharedReg1221_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1221_out;
   MUX_Add30_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1156_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1221_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1002_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg991_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1221_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1059_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1002_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1000_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg599_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay96No2_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg642_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1227_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg425_out_to_MUX_Add30_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_2_impl_1_out);

   Delay1No221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_2_impl_1_out,
                 Y => Delay1No221_out);

Delay1No222_out_to_Add30_3_impl_parent_implementedSystem_port_0_cast <= Delay1No222_out;
Delay1No223_out_to_Add30_3_impl_parent_implementedSystem_port_1_cast <= Delay1No223_out;
   Add30_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_3_impl_out,
                 X => Delay1No222_out_to_Add30_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No223_out_to_Add30_3_impl_parent_implementedSystem_port_1_cast);

Delay24No2_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_1_cast <= Delay24No2_out;
Delay73No8_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_2_cast <= Delay73No8_out;
SharedReg751_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg751_out;
SharedReg551_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg551_out;
SharedReg690_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg690_out;
SharedReg608_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg608_out;
SharedReg761_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg761_out;
SharedReg609_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg609_out;
SharedReg605_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg605_out;
SharedReg561_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg561_out;
SharedReg656_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg656_out;
SharedReg1160_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1160_out;
SharedReg379_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg379_out;
   MUX_Add30_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay24No2_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay73No8_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg656_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1160_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg379_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg751_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg551_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg690_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg608_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg761_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg609_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg605_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg561_out_to_MUX_Add30_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_3_impl_0_out);

   Delay1No222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_3_impl_0_out,
                 Y => Delay1No222_out);

SharedReg1229_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1229_out;
SharedReg1227_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1227_out;
SharedReg1163_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1163_out;
SharedReg1227_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1227_out;
SharedReg423_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg423_out;
SharedReg1232_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1232_out;
SharedReg1037_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1037_out;
SharedReg654_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg654_out;
Delay96No3_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_9_cast <= Delay96No3_out;
SharedReg755_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg755_out;
SharedReg1233_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1233_out;
SharedReg1002_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1002_out;
SharedReg598_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg598_out;
   MUX_Add30_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1229_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1227_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1233_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1002_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg598_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1163_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1227_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg423_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1232_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1037_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg654_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay96No3_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg755_out_to_MUX_Add30_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_3_impl_1_out);

   Delay1No223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_3_impl_1_out,
                 Y => Delay1No223_out);

Delay1No224_out_to_Add30_4_impl_parent_implementedSystem_port_0_cast <= Delay1No224_out;
Delay1No225_out_to_Add30_4_impl_parent_implementedSystem_port_1_cast <= Delay1No225_out;
   Add30_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_4_impl_out,
                 X => Delay1No224_out_to_Add30_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No225_out_to_Add30_4_impl_parent_implementedSystem_port_1_cast);

SharedReg1167_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1167_out;
SharedReg437_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg437_out;
Delay60No3_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_3_cast <= Delay60No3_out;
SharedReg808_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg808_out;
SharedReg485_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg485_out;
Delay104No3_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_6_cast <= Delay104No3_out;
Delay88No10_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_7_cast <= Delay88No10_out;
SharedReg1182_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1182_out;
Delay69No10_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_9_cast <= Delay69No10_out;
SharedReg445_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg445_out;
SharedReg1198_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1198_out;
SharedReg571_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg571_out;
SharedReg436_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg436_out;
   MUX_Add30_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1167_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg437_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1198_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg571_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg436_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay60No3_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg808_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg485_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay104No3_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay88No10_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1182_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay69No10_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg445_out_to_MUX_Add30_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_4_impl_0_out);

   Delay1No224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_4_impl_0_out,
                 Y => Delay1No224_out);

SharedReg1127_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1127_out;
SharedReg1127_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1127_out;
SharedReg1127_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1127_out;
SharedReg957_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg957_out;
SharedReg1094_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1094_out;
SharedReg1234_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1234_out;
SharedReg1097_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1097_out;
SharedReg1236_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1236_out;
SharedReg1097_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1097_out;
SharedReg968_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg968_out;
SharedReg1236_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1236_out;
SharedReg762_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg762_out;
SharedReg1091_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1091_out;
   MUX_Add30_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1127_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1127_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1236_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg762_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1091_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1127_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg957_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1094_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1234_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1097_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1236_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1097_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg968_out_to_MUX_Add30_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_4_impl_1_out);

   Delay1No225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_4_impl_1_out,
                 Y => Delay1No225_out);

Delay1No226_out_to_Add30_5_impl_parent_implementedSystem_port_0_cast <= Delay1No226_out;
Delay1No227_out_to_Add30_5_impl_parent_implementedSystem_port_1_cast <= Delay1No227_out;
   Add30_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add30_5_impl_out,
                 X => Delay1No226_out_to_Add30_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No227_out_to_Add30_5_impl_parent_implementedSystem_port_1_cast);

Delay5No16_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_1_cast <= Delay5No16_out;
SharedReg528_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg528_out;
SharedReg526_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg526_out;
SharedReg1211_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1211_out;
Delay60No4_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_5_cast <= Delay60No4_out;
Delay89No10_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_6_cast <= Delay89No10_out;
SharedReg1180_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1180_out;
SharedReg1175_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1175_out;
Delay104No11_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_9_cast <= Delay104No11_out;
SharedReg1262_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1262_out;
SharedReg670_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg670_out;
SharedReg672_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg672_out;
SharedReg448_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg448_out;
   MUX_Add30_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No16_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg528_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg670_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg672_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg448_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg526_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1211_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay60No4_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay89No10_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1180_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1175_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay104No11_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1262_out_to_MUX_Add30_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_5_impl_0_out);

   Delay1No226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_5_impl_0_out,
                 Y => Delay1No226_out);

SharedReg487_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg487_out;
SharedReg669_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg669_out;
Delay70No5_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_3_cast <= Delay70No5_out;
SharedReg1248_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1248_out;
SharedReg968_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg968_out;
SharedReg1071_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1071_out;
SharedReg1115_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1115_out;
SharedReg1115_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1115_out;
SharedReg1247_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1247_out;
SharedReg1104_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1104_out;
SharedReg398_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg398_out;
SharedReg1244_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1244_out;
SharedReg968_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg968_out;
   MUX_Add30_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg487_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg669_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg398_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1244_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg968_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay70No5_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1248_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg968_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1071_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1115_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1115_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1247_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1104_out_to_MUX_Add30_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add30_5_impl_1_out);

   Delay1No227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add30_5_impl_1_out,
                 Y => Delay1No227_out);

Delay1No228_out_to_Add110_1_impl_parent_implementedSystem_port_0_cast <= Delay1No228_out;
Delay1No229_out_to_Add110_1_impl_parent_implementedSystem_port_1_cast <= Delay1No229_out;
   Add110_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add110_1_impl_out,
                 X => Delay1No228_out_to_Add110_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No229_out_to_Add110_1_impl_parent_implementedSystem_port_1_cast);

SharedReg627_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg627_out;
SharedReg592_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg592_out;
SharedReg744_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg744_out;
SharedReg593_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg593_out;
Delay55No6_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_5_cast <= Delay55No6_out;
Delay5No12_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_6_cast <= Delay5No12_out;
SharedReg410_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg410_out;
Delay19No13_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_8_cast <= Delay19No13_out;
SharedReg635_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg635_out;
SharedReg540_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg540_out;
SharedReg371_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg371_out;
Delay69No12_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_12_cast <= Delay69No12_out;
SharedReg494_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg494_out;
   MUX_Add110_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg627_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg592_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg371_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay69No12_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg494_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg744_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg593_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay55No6_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay5No12_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg410_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay19No13_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg635_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg540_out_to_MUX_Add110_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add110_1_impl_0_out);

   Delay1No228_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_1_impl_0_out,
                 Y => Delay1No228_out);

SharedReg404_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg404_out;
SharedReg1220_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1220_out;
SharedReg987_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg987_out;
SharedReg591_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg591_out;
SharedReg991_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg991_out;
SharedReg363_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg363_out;
Delay70No1_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_7_cast <= Delay70No1_out;
SharedReg943_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg943_out;
SharedReg887_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg887_out;
SharedReg592_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg592_out;
SharedReg590_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg590_out;
SharedReg1082_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1082_out;
SharedReg359_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg359_out;
   MUX_Add110_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg404_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1220_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg590_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1082_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg359_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg987_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg591_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg991_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg363_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay70No1_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg943_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg887_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg592_out_to_MUX_Add110_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add110_1_impl_1_out);

   Delay1No229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_1_impl_1_out,
                 Y => Delay1No229_out);

Delay1No230_out_to_Add110_2_impl_parent_implementedSystem_port_0_cast <= Delay1No230_out;
Delay1No231_out_to_Add110_2_impl_parent_implementedSystem_port_1_cast <= Delay1No231_out;
   Add110_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add110_2_impl_out,
                 X => Delay1No230_out_to_Add110_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No231_out_to_Add110_2_impl_parent_implementedSystem_port_1_cast);

SharedReg415_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg415_out;
SharedReg500_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg500_out;
SharedReg634_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg634_out;
SharedReg600_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg600_out;
SharedReg375_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg375_out;
SharedReg1158_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1158_out;
Delay55No7_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_7_cast <= Delay55No7_out;
Delay5No13_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_8_cast <= Delay5No13_out;
SharedReg420_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg420_out;
SharedReg1166_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1166_out;
SharedReg747_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg747_out;
SharedReg1153_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1153_out;
SharedReg880_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg880_out;
   MUX_Add110_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg415_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg500_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg747_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1153_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg880_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg634_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg600_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg375_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1158_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay55No7_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay5No13_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg420_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1166_out_to_MUX_Add110_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add110_2_impl_0_out);

   Delay1No230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_2_impl_0_out,
                 Y => Delay1No230_out);

SharedReg594_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg594_out;
SharedReg458_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg458_out;
SharedReg413_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg413_out;
SharedReg1226_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1226_out;
SharedReg1218_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1218_out;
SharedReg1002_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1002_out;
SharedReg1002_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1002_out;
SharedReg418_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg418_out;
Delay70No2_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_9_cast <= Delay70No2_out;
SharedReg1091_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1091_out;
SharedReg893_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg893_out;
SharedReg371_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg371_out;
SharedReg1137_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1137_out;
   MUX_Add110_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg594_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg458_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg893_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg371_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1137_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg413_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1226_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1218_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1002_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1002_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg418_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay70No2_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1091_out_to_MUX_Add110_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add110_2_impl_1_out);

   Delay1No231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_2_impl_1_out,
                 Y => Delay1No231_out);

Delay1No232_out_to_Add110_3_impl_parent_implementedSystem_port_0_cast <= Delay1No232_out;
Delay1No233_out_to_Add110_3_impl_parent_implementedSystem_port_1_cast <= Delay1No233_out;
   Add110_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add110_3_impl_out,
                 X => Delay1No232_out_to_Add110_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No233_out_to_Add110_3_impl_parent_implementedSystem_port_1_cast);

SharedReg892_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg892_out;
SharedReg888_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg888_out;
SharedReg469_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg469_out;
SharedReg505_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg505_out;
SharedReg699_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg699_out;
SharedReg385_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg385_out;
SharedReg383_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg383_out;
SharedReg1165_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1165_out;
Delay55No8_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_9_cast <= Delay55No8_out;
Delay5No14_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_10_cast <= Delay5No14_out;
SharedReg559_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg559_out;
Delay88No2_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_12_cast <= Delay88No2_out;
SharedReg745_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg745_out;
   MUX_Add110_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg892_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg888_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg559_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay88No2_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg745_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg469_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg505_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg699_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg385_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg383_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1165_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay55No8_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay5No14_out_to_MUX_Add110_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add110_3_impl_0_out);

   Delay1No232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_3_impl_0_out,
                 Y => Delay1No232_out);

SharedReg1059_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1059_out;
SharedReg1059_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1059_out;
SharedReg602_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg602_out;
SharedReg465_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg465_out;
SharedReg1021_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1021_out;
SharedReg1127_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1127_out;
SharedReg1224_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1224_out;
SharedReg1127_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1127_out;
SharedReg1127_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1127_out;
SharedReg511_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg511_out;
Delay70No3_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_11_cast <= Delay70No3_out;
SharedReg1225_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1225_out;
SharedReg934_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg934_out;
   MUX_Add110_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1059_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1059_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay70No3_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1225_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg934_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg602_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg465_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1021_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1127_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1224_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1127_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1127_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg511_out_to_MUX_Add110_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add110_3_impl_1_out);

   Delay1No233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_3_impl_1_out,
                 Y => Delay1No233_out);

Delay1No234_out_to_Add110_4_impl_parent_implementedSystem_port_0_cast <= Delay1No234_out;
Delay1No235_out_to_Add110_4_impl_parent_implementedSystem_port_1_cast <= Delay1No235_out;
   Add110_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add110_4_impl_out,
                 X => Delay1No234_out_to_Add110_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No235_out_to_Add110_4_impl_parent_implementedSystem_port_1_cast);

SharedReg446_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg446_out;
SharedReg763_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg763_out;
SharedReg566_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg566_out;
SharedReg1191_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1191_out;
SharedReg906_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg906_out;
SharedReg1168_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1168_out;
SharedReg616_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg616_out;
SharedReg567_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg567_out;
SharedReg862_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg862_out;
Delay88No11_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_10_cast <= Delay88No11_out;
SharedReg672_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg672_out;
SharedReg568_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg568_out;
SharedReg568_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg568_out;
   MUX_Add110_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg446_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg763_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg672_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg568_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg568_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg566_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1191_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg906_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1168_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg616_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg567_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg862_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay88No11_out_to_MUX_Add110_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add110_4_impl_0_out);

   Delay1No234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_4_impl_0_out,
                 Y => Delay1No234_out);

SharedReg1070_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1070_out;
SharedReg907_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg907_out;
SharedReg764_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg764_out;
SharedReg611_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg611_out;
SharedReg965_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg965_out;
SharedReg965_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg965_out;
SharedReg613_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg613_out;
SharedReg481_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg481_out;
Delay67No4_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_9_cast <= Delay67No4_out;
SharedReg971_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg971_out;
SharedReg1244_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1244_out;
SharedReg1011_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1011_out;
Delay70No4_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_13_cast <= Delay70No4_out;
   MUX_Add110_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1070_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg907_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1244_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1011_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay70No4_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg764_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg611_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg965_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg965_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg613_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg481_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay67No4_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg971_out_to_MUX_Add110_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add110_4_impl_1_out);

   Delay1No235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add110_4_impl_1_out,
                 Y => Delay1No235_out);

Delay1No236_out_to_Add101_2_impl_parent_implementedSystem_port_0_cast <= Delay1No236_out;
Delay1No237_out_to_Add101_2_impl_parent_implementedSystem_port_1_cast <= Delay1No237_out;
   Add101_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add101_2_impl_out,
                 X => Delay1No236_out_to_Add101_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No237_out_to_Add101_2_impl_parent_implementedSystem_port_1_cast);

SharedReg468_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg468_out;
Delay104No1_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_2_cast <= Delay104No1_out;
Delay88No8_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_3_cast <= Delay88No8_out;
SharedReg799_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg799_out;
SharedReg507_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg507_out;
SharedReg1162_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1162_out;
SharedReg692_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg692_out;
SharedReg420_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg420_out;
SharedReg603_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg603_out;
Delay5No8_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_10_cast <= Delay5No8_out;
SharedReg1163_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1163_out;
SharedReg550_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg550_out;
Delay104No7_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_13_cast <= Delay104No7_out;
   MUX_Add101_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg468_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay104No1_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1163_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg550_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay104No7_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay88No8_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg799_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg507_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1162_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg692_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg420_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg603_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay5No8_out_to_MUX_Add101_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add101_2_impl_0_out);

   Delay1No236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_2_impl_0_out,
                 Y => Delay1No236_out);

SharedReg933_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg933_out;
SharedReg1222_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1222_out;
SharedReg1021_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1021_out;
SharedReg1224_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1224_out;
SharedReg1226_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1226_out;
SharedReg1091_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1091_out;
SharedReg754_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg754_out;
SharedReg1002_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1002_out;
SharedReg1225_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1225_out;
SharedReg471_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg471_out;
SharedReg1017_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1017_out;
SharedReg749_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg749_out;
SharedReg1223_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1223_out;
   MUX_Add101_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg933_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1222_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1017_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg749_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1223_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1021_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1224_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1226_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1091_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg754_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1002_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1225_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg471_out_to_MUX_Add101_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add101_2_impl_1_out);

   Delay1No237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_2_impl_1_out,
                 Y => Delay1No237_out);

Delay1No238_out_to_Add101_3_impl_parent_implementedSystem_port_0_cast <= Delay1No238_out;
Delay1No239_out_to_Add101_3_impl_parent_implementedSystem_port_1_cast <= Delay1No239_out;
   Add101_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add101_3_impl_out,
                 X => Delay1No238_out_to_Add101_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No239_out_to_Add101_3_impl_parent_implementedSystem_port_1_cast);

SharedReg557_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg557_out;
SharedReg386_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg386_out;
SharedReg563_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg563_out;
Delay73No9_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_4_cast <= Delay73No9_out;
Delay76No3_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_5_cast <= Delay76No3_out;
SharedReg558_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg558_out;
SharedReg700_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg700_out;
SharedReg664_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg664_out;
SharedReg768_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg768_out;
SharedReg665_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg665_out;
SharedReg610_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg610_out;
Delay5No9_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_12_cast <= Delay5No9_out;
SharedReg756_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg756_out;
   MUX_Add101_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg557_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg386_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg610_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay5No9_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg756_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg563_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay73No9_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay76No3_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg558_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg700_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg664_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg768_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg665_out_to_MUX_Add101_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add101_3_impl_0_out);

   Delay1No238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_3_impl_0_out,
                 Y => Delay1No238_out);

SharedReg757_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg757_out;
SharedReg606_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg606_out;
SharedReg1235_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1235_out;
SharedReg1233_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1233_out;
Delay6No3_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_5_cast <= Delay6No3_out;
SharedReg474_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg474_out;
SharedReg476_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg476_out;
SharedReg1238_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1238_out;
SharedReg1016_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1016_out;
SharedReg711_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg711_out;
Delay96No4_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_11_cast <= Delay96No4_out;
SharedReg479_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg479_out;
SharedReg901_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg901_out;
   MUX_Add101_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg757_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg606_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay96No4_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg479_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg901_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1235_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1233_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay6No3_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg474_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg476_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1238_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1016_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg711_out_to_MUX_Add101_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add101_3_impl_1_out);

   Delay1No239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_3_impl_1_out,
                 Y => Delay1No239_out);

Delay1No240_out_to_Add101_5_impl_parent_implementedSystem_port_0_cast <= Delay1No240_out;
Delay1No241_out_to_Add101_5_impl_parent_implementedSystem_port_1_cast <= Delay1No241_out;
   Add101_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add101_5_impl_out,
                 X => Delay1No240_out_to_Add101_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No241_out_to_Add101_5_impl_parent_implementedSystem_port_1_cast);

SharedReg573_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg573_out;
SharedReg526_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg526_out;
SharedReg823_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg823_out;
Delay5No5_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_4_cast <= Delay5No5_out;
SharedReg719_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg719_out;
SharedReg487_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg487_out;
SharedReg1200_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1200_out;
SharedReg675_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg675_out;
SharedReg923_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg923_out;
SharedReg1210_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1210_out;
SharedReg719_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg719_out;
Delay69No11_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_12_cast <= Delay69No11_out;
SharedReg772_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg772_out;
   MUX_Add101_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg573_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg526_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg719_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay69No11_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg772_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg823_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay5No5_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg719_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg487_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1200_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg675_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg923_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1210_out_to_MUX_Add101_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add101_5_impl_0_out);

   Delay1No240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_5_impl_0_out,
                 Y => Delay1No240_out);

Delay96No5_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_1_cast <= Delay96No5_out;
SharedReg1070_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1070_out;
SharedReg1245_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1245_out;
SharedReg1200_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1200_out;
SharedReg871_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg871_out;
SharedReg720_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg720_out;
SharedReg525_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg525_out;
SharedReg1247_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1247_out;
SharedReg1045_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1045_out;
SharedReg1248_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1248_out;
SharedReg1245_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1245_out;
SharedReg1108_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1108_out;
SharedReg771_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg771_out;
   MUX_Add101_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay96No5_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1070_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1245_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1108_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg771_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1245_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1200_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg871_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg720_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg525_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1247_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1045_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1248_out_to_MUX_Add101_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add101_5_impl_1_out);

   Delay1No241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add101_5_impl_1_out,
                 Y => Delay1No241_out);

Delay1No242_out_to_Add111_1_impl_parent_implementedSystem_port_0_cast <= Delay1No242_out;
Delay1No243_out_to_Add111_1_impl_parent_implementedSystem_port_1_cast <= Delay1No243_out;
   Add111_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add111_1_impl_out,
                 X => Delay1No242_out_to_Add111_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No243_out_to_Add111_1_impl_parent_implementedSystem_port_1_cast);

Delay88No7_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_1_cast <= Delay88No7_out;
Delay76No7_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_2_cast <= Delay76No7_out;
SharedReg689_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg689_out;
SharedReg1159_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1159_out;
SharedReg686_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg686_out;
SharedReg365_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg365_out;
SharedReg595_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg595_out;
Delay5No7_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_8_cast <= Delay5No7_out;
SharedReg889_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg889_out;
SharedReg1153_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1153_out;
SharedReg890_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg890_out;
Delay24No1_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_12_cast <= Delay24No1_out;
Delay104No_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_13_cast <= Delay104No_out;
   MUX_Add111_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay88No7_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay76No7_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg890_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay24No1_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay104No_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg689_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1159_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg686_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg365_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg595_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay5No7_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg889_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1153_out_to_MUX_Add111_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add111_1_impl_0_out);

   Delay1No242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_1_impl_0_out,
                 Y => Delay1No242_out);

SharedReg937_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg937_out;
SharedReg1218_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1218_out;
SharedReg1062_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1062_out;
SharedReg943_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg943_out;
SharedReg744_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg744_out;
SharedReg991_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg991_out;
SharedReg1219_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1219_out;
SharedReg371_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg371_out;
SharedReg933_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg933_out;
SharedReg991_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg991_out;
SharedReg991_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg991_out;
SharedReg1223_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1223_out;
SharedReg1216_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1216_out;
   MUX_Add111_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg937_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1218_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg991_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1223_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1216_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1062_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg943_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg744_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg991_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1219_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg371_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg933_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg991_out_to_MUX_Add111_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add111_1_impl_1_out);

   Delay1No243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_1_impl_1_out,
                 Y => Delay1No243_out);

Delay1No244_out_to_Add111_4_impl_parent_implementedSystem_port_0_cast <= Delay1No244_out;
Delay1No245_out_to_Add111_4_impl_parent_implementedSystem_port_1_cast <= Delay1No245_out;
   Add111_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add111_4_impl_out,
                 X => Delay1No244_out_to_Add111_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No245_out_to_Add111_4_impl_parent_implementedSystem_port_1_cast);

Delay5No4_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_1_cast <= Delay5No4_out;
SharedReg442_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg442_out;
Delay88No4_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_3_cast <= Delay88No4_out;
Delay14No4_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_4_cast <= Delay14No4_out;
SharedReg615_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg615_out;
Delay73No10_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_6_cast <= Delay73No10_out;
SharedReg766_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg766_out;
SharedReg611_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg611_out;
SharedReg447_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg447_out;
SharedReg579_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg579_out;
SharedReg580_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg580_out;
SharedReg1196_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1196_out;
SharedReg714_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg714_out;
   MUX_Add111_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No4_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg442_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg580_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1196_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg714_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay88No4_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay14No4_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg615_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay73No10_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg766_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg611_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg447_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg579_out_to_MUX_Add111_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add111_4_impl_0_out);

   Delay1No244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_4_impl_0_out,
                 Y => Delay1No244_out);

SharedReg394_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg394_out;
SharedReg965_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg965_out;
SharedReg1237_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1237_out;
SharedReg716_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg716_out;
SharedReg1241_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1241_out;
SharedReg1239_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1239_out;
SharedReg1176_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1176_out;
SharedReg1239_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1239_out;
SharedReg1115_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1115_out;
SharedReg576_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg576_out;
SharedReg1104_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1104_out;
SharedReg968_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg968_out;
SharedReg1239_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1239_out;
   MUX_Add111_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg394_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg965_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1104_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg968_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1239_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1237_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg716_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1241_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1239_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1176_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1239_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1115_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg576_out_to_MUX_Add111_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add111_4_impl_1_out);

   Delay1No245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add111_4_impl_1_out,
                 Y => Delay1No245_out);

Delay1No246_out_to_Add141_0_impl_parent_implementedSystem_port_0_cast <= Delay1No246_out;
Delay1No247_out_to_Add141_0_impl_parent_implementedSystem_port_1_cast <= Delay1No247_out;
   Add141_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add141_0_impl_out,
                 X => Delay1No246_out_to_Add141_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No247_out_to_Add141_0_impl_parent_implementedSystem_port_1_cast);

SharedReg496_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg496_out;
SharedReg1150_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1150_out;
SharedReg678_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg678_out;
SharedReg356_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg356_out;
SharedReg631_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg631_out;
Delay5No_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_6_cast <= Delay5No_out;
SharedReg1148_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1148_out;
Delay88No_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_8_cast <= Delay88No_out;
SharedReg412_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg412_out;
SharedReg1148_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1148_out;
Delay104No6_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_11_cast <= Delay104No6_out;
SharedReg406_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg406_out;
SharedReg407_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg407_out;
   MUX_Add141_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg496_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1150_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay104No6_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg406_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg407_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg678_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg356_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg631_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay5No_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1148_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay88No_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg412_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1148_out_to_MUX_Add141_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add141_0_impl_0_out);

   Delay1No246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add141_0_impl_0_out,
                 Y => Delay1No246_out);

SharedReg1214_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1214_out;
SharedReg1082_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1082_out;
SharedReg732_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg732_out;
SharedReg1082_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1082_out;
SharedReg1215_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1215_out;
SharedReg879_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg879_out;
SharedReg1137_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1137_out;
SharedReg1213_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1213_out;
SharedReg632_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg632_out;
SharedReg363_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg363_out;
SharedReg1217_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1217_out;
SharedReg453_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg453_out;
SharedReg1082_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1082_out;
   MUX_Add141_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1214_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1082_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1217_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg453_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1082_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg732_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1082_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1215_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg879_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1137_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1213_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg632_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg363_out_to_MUX_Add141_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add141_0_impl_1_out);

   Delay1No247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add141_0_impl_1_out,
                 Y => Delay1No247_out);

Delay1No248_out_to_Add141_2_impl_parent_implementedSystem_port_0_cast <= Delay1No248_out;
Delay1No249_out_to_Add141_2_impl_parent_implementedSystem_port_1_cast <= Delay1No249_out;
   Add141_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add141_2_impl_out,
                 X => Delay1No248_out_to_Add141_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No249_out_to_Add141_2_impl_parent_implementedSystem_port_1_cast);

SharedReg1160_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1160_out;
Delay104No8_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_2_cast <= Delay104No8_out;
SharedReg477_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg477_out;
Delay104No2_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_4_cast <= Delay104No2_out;
SharedReg475_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg475_out;
SharedReg478_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg478_out;
SharedReg513_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg513_out;
SharedReg388_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg388_out;
SharedReg757_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg757_out;
SharedReg473_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg473_out;
SharedReg655_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg655_out;
SharedReg1173_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1173_out;
SharedReg430_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg430_out;
   MUX_Add141_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1160_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay104No8_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg655_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1173_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg430_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg477_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay104No2_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg475_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg478_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg513_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg388_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg757_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg473_out_to_MUX_Add141_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add141_2_impl_0_out);

   Delay1No248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add141_2_impl_0_out,
                 Y => Delay1No248_out);

SharedReg379_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg379_out;
SharedReg1229_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1229_out;
SharedReg943_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg943_out;
SharedReg1228_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1228_out;
SharedReg1127_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1127_out;
SharedReg1094_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1094_out;
SharedReg1232_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1232_out;
SharedReg1094_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1094_out;
SharedReg761_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg761_out;
SharedReg1028_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1028_out;
SharedReg1231_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1231_out;
SharedReg1094_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1094_out;
SharedReg649_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg649_out;
   MUX_Add141_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg379_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1229_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1231_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1094_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg649_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg943_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1228_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1127_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1094_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1232_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1094_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg761_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1028_out_to_MUX_Add141_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add141_2_impl_1_out);

   Delay1No249_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add141_2_impl_1_out,
                 Y => Delay1No249_out);

Delay1No250_out_to_Add141_3_impl_parent_implementedSystem_port_0_cast <= Delay1No250_out;
Delay1No251_out_to_Add141_3_impl_parent_implementedSystem_port_1_cast <= Delay1No251_out;
   Add141_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add141_3_impl_out,
                 X => Delay1No250_out_to_Add141_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No251_out_to_Add141_3_impl_parent_implementedSystem_port_1_cast);

Delay88No3_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_1_cast <= Delay88No3_out;
SharedReg440_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg440_out;
SharedReg1167_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1167_out;
Delay104No9_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_4_cast <= Delay104No9_out;
SharedReg759_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg759_out;
SharedReg606_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg606_out;
SharedReg483_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg483_out;
SharedReg617_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg617_out;
SharedReg569_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg569_out;
SharedReg395_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg395_out;
SharedReg811_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg811_out;
Delay5No15_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_12_cast <= Delay5No15_out;
SharedReg479_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg479_out;
   MUX_Add141_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay88No3_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg440_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg811_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay5No15_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg479_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1167_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay104No9_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg759_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg606_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg483_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg617_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg569_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg395_out_to_MUX_Add141_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add141_3_impl_0_out);

   Delay1No250_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add141_3_impl_0_out,
                 Y => Delay1No250_out);

SharedReg1231_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1231_out;
SharedReg658_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg658_out;
SharedReg386_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg386_out;
SharedReg1235_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1235_out;
SharedReg1170_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1170_out;
SharedReg1233_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1233_out;
SharedReg965_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg965_out;
SharedReg1070_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1070_out;
SharedReg1238_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1238_out;
SharedReg1115_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1115_out;
SharedReg817_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg817_out;
SharedReg517_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg517_out;
SharedReg1127_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1127_out;
   MUX_Add141_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1231_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg658_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg817_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg517_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1127_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg386_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1235_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1170_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1233_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg965_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1070_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1238_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1115_out_to_MUX_Add141_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add141_3_impl_1_out);

   Delay1No251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add141_3_impl_1_out,
                 Y => Delay1No251_out);

Delay1No252_out_to_Add141_5_impl_parent_implementedSystem_port_0_cast <= Delay1No252_out;
Delay1No253_out_to_Add141_5_impl_parent_implementedSystem_port_1_cast <= Delay1No253_out;
   Add141_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add141_5_impl_out,
                 X => Delay1No252_out_to_Add141_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No253_out_to_Add141_5_impl_parent_implementedSystem_port_1_cast);

Delay5No11_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_1_cast <= Delay5No11_out;
Delay88No5_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_2_cast <= Delay88No5_out;
Delay104No5_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_3_cast <= Delay104No5_out;
SharedReg774_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg774_out;
SharedReg819_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg819_out;
SharedReg1209_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1209_out;
SharedReg874_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg874_out;
SharedReg1259_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1259_out;
SharedReg1260_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1260_out;
SharedReg1207_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1207_out;
SharedReg1200_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1200_out;
   MUX_Add141_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_11_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No11_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay88No5_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1200_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_2 => Delay104No5_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg774_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg819_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1209_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg874_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1259_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1260_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1207_out_to_MUX_Add141_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add141_5_impl_0_LUT_out,
                 oMux => MUX_Add141_5_impl_0_out);

   Delay1No252_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add141_5_impl_0_out,
                 Y => Delay1No252_out);

SharedReg578_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg578_out;
SharedReg724_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg724_out;
SharedReg825_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg825_out;
SharedReg1243_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1243_out;
SharedReg1246_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1246_out;
SharedReg1243_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1243_out;
SharedReg1104_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1104_out;
SharedReg1248_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1248_out;
SharedReg1044_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1044_out;
SharedReg1207_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1207_out;
SharedReg1207_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1207_out;
   MUX_Add141_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_11_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg578_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg724_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1207_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_2 => SharedReg825_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1243_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1246_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1243_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1104_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1248_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1044_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1207_out_to_MUX_Add141_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add141_5_impl_1_LUT_out,
                 oMux => MUX_Add141_5_impl_1_out);

   Delay1No253_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add141_5_impl_1_out,
                 Y => Delay1No253_out);

Delay1No254_out_to_Add151_5_impl_parent_implementedSystem_port_0_cast <= Delay1No254_out;
Delay1No255_out_to_Add151_5_impl_parent_implementedSystem_port_1_cast <= Delay1No255_out;
   Add151_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add151_5_impl_out,
                 X => Delay1No254_out_to_Add151_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No255_out_to_Add151_5_impl_parent_implementedSystem_port_1_cast);

Delay5No10_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_1_cast <= Delay5No10_out;
SharedReg396_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg396_out;
SharedReg1174_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1174_out;
SharedReg397_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg397_out;
SharedReg1191_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1191_out;
SharedReg818_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg818_out;
SharedReg449_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg449_out;
SharedReg818_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg818_out;
Delay73No11_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_9_cast <= Delay73No11_out;
SharedReg722_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg722_out;
SharedReg922_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg922_out;
Delay59No5_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_12_cast <= Delay59No5_out;
SharedReg667_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg667_out;
   MUX_Add151_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No10_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg396_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg922_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay59No5_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg667_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1174_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg397_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1191_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg818_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg449_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg818_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay73No11_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg722_out_to_MUX_Add151_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add151_5_impl_0_out);

   Delay1No254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add151_5_impl_0_out,
                 Y => Delay1No254_out);

SharedReg442_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg442_out;
SharedReg1094_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1094_out;
SharedReg965_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg965_out;
SharedReg1070_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1070_out;
SharedReg394_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg394_out;
SharedReg1241_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1241_out;
SharedReg1070_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1070_out;
SharedReg1240_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1240_out;
SharedReg1245_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1245_out;
SharedReg1185_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1185_out;
SharedReg1242_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1242_out;
SharedReg1054_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1054_out;
SharedReg1237_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1237_out;
   MUX_Add151_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg442_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1094_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1242_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1054_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1237_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg965_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1070_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg394_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1241_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1070_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1240_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1245_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1185_out_to_MUX_Add151_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add151_5_impl_1_out);

   Delay1No255_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add151_5_impl_1_out,
                 Y => Delay1No255_out);

Delay1No256_out_to_Add21_3_impl_parent_implementedSystem_port_0_cast <= Delay1No256_out;
Delay1No257_out_to_Add21_3_impl_parent_implementedSystem_port_1_cast <= Delay1No257_out;
   Add21_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add21_3_impl_out,
                 X => Delay1No256_out_to_Add21_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No257_out_to_Add21_3_impl_parent_implementedSystem_port_1_cast);

SharedReg850_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg850_out;
Delay89No8_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_2_cast <= Delay89No8_out;
Delay15No26_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_3_cast <= Delay15No26_out;
SharedReg894_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg894_out;
Delay88No9_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_5_cast <= Delay88No9_out;
Delay76No9_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_6_cast <= Delay76No9_out;
SharedReg708_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg708_out;
SharedReg482_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg482_out;
SharedReg392_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg392_out;
SharedReg391_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg391_out;
SharedReg484_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg484_out;
Delay5No3_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_12_cast <= Delay5No3_out;
SharedReg428_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg428_out;
   MUX_Add21_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg850_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay89No8_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg484_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay5No3_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg428_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay15No26_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg894_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay88No9_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay76No9_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg708_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg482_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg392_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg391_out_to_MUX_Add21_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add21_3_impl_0_out);

   Delay1No256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add21_3_impl_0_out,
                 Y => Delay1No256_out);

SharedReg1002_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1002_out;
SharedReg944_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg944_out;
SharedReg1017_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1017_out;
SharedReg956_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg956_out;
SharedReg1093_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1093_out;
SharedReg1230_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1230_out;
SharedReg1093_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1093_out;
SharedReg965_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg965_out;
SharedReg1230_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1230_out;
SharedReg1011_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1011_out;
SharedReg1011_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1011_out;
SharedReg433_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg433_out;
SharedReg1002_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1002_out;
   MUX_Add21_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1002_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg944_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1011_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg433_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1002_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1017_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg956_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1093_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1230_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1093_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg965_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1230_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1011_out_to_MUX_Add21_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add21_3_impl_1_out);

   Delay1No257_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add21_3_impl_1_out,
                 Y => Delay1No257_out);

Delay1No258_out_to_Add23_0_impl_parent_implementedSystem_port_0_cast <= Delay1No258_out;
Delay1No259_out_to_Add23_0_impl_parent_implementedSystem_port_1_cast <= Delay1No259_out;
   Add23_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add23_0_impl_out,
                 X => Delay1No258_out_to_Add23_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No259_out_to_Add23_0_impl_parent_implementedSystem_port_1_cast);

SharedReg683_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg683_out;
SharedReg884_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg884_out;
SharedReg883_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg883_out;
SharedReg1152_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1152_out;
SharedReg587_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg587_out;
Delay5No6_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_6_cast <= Delay5No6_out;
SharedReg829_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg829_out;
SharedReg827_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg827_out;
SharedReg882_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg882_out;
Delay60No_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_10_cast <= Delay60No_out;
SharedReg734_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg734_out;
SharedReg586_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg586_out;
SharedReg733_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg733_out;
   MUX_Add23_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg683_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg884_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg734_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg586_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg733_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg883_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1152_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg587_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay5No6_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg829_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg827_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg882_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => Delay60No_out_to_MUX_Add23_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add23_0_impl_0_out);

   Delay1No258_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add23_0_impl_0_out,
                 Y => Delay1No258_out);

SharedReg1086_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1086_out;
SharedReg1137_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1137_out;
SharedReg1212_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1212_out;
SharedReg933_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg933_out;
SharedReg1213_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1213_out;
SharedReg1148_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1148_out;
SharedReg1082_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1082_out;
SharedReg1137_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1137_out;
SharedReg1137_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1137_out;
SharedReg977_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg977_out;
SharedReg1083_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1083_out;
SharedReg1151_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1151_out;
SharedReg1212_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1212_out;
   MUX_Add23_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1086_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1137_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1083_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1151_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1212_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1212_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg933_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1213_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1148_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1082_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1137_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1137_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg977_out_to_MUX_Add23_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Add23_0_impl_1_out);

   Delay1No259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add23_0_impl_1_out,
                 Y => Delay1No259_out);

Delay1No260_out_to_Product312_0_impl_parent_implementedSystem_port_0_cast <= Delay1No260_out;
Delay1No261_out_to_Product312_0_impl_parent_implementedSystem_port_1_cast <= Delay1No261_out;
   Product312_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product312_0_impl_out,
                 X => Delay1No260_out_to_Product312_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No261_out_to_Product312_0_impl_parent_implementedSystem_port_1_cast);

SharedReg6_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg6_out;
Delay1No338_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_2_cast <= Delay1No338_out;
SharedReg880_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg880_out;
SharedReg778_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg778_out;
SharedReg400_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg400_out;
SharedReg726_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg726_out;
SharedReg681_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg681_out;
SharedReg726_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg726_out;
SharedReg881_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg881_out;
SharedReg241_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg241_out;
SharedReg977_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg977_out;
SharedReg828_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg828_out;
SharedReg4_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg4_out;
   MUX_Product312_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg6_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No338_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg977_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg828_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg4_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg880_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg778_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg400_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg726_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg681_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg726_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg881_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg241_out_to_MUX_Product312_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product312_0_impl_0_out);

   Delay1No260_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product312_0_impl_0_out,
                 Y => Delay1No260_out);

SharedReg181_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg181_out;
SharedReg1263_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1263_out;
SharedReg1314_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1314_out;
SharedReg1288_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1288_out;
SharedReg242_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg242_out;
SharedReg1278_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1278_out;
SharedReg1279_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1279_out;
SharedReg1292_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1292_out;
SharedReg1281_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1281_out;
SharedReg177_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg177_out;
SharedReg1137_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1137_out;
SharedReg1272_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1272_out;
SharedReg978_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg978_out;
   MUX_Product312_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg181_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1263_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1137_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1272_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg978_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1314_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1288_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg242_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1278_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1279_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1292_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1281_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg177_out_to_MUX_Product312_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product312_0_impl_1_out);

   Delay1No261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product312_0_impl_1_out,
                 Y => Delay1No261_out);

Delay1No262_out_to_Product312_1_impl_parent_implementedSystem_port_0_cast <= Delay1No262_out;
Delay1No263_out_to_Product312_1_impl_parent_implementedSystem_port_1_cast <= Delay1No263_out;
   Product312_1_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product312_1_impl_out,
                 X => Delay1No262_out_to_Product312_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No263_out_to_Product312_1_impl_parent_implementedSystem_port_1_cast);

SharedReg835_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg835_out;
SharedReg424_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg424_out;
SharedReg17_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg17_out;
Delay1No333_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_4_cast <= Delay1No333_out;
SharedReg936_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg936_out;
SharedReg790_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg790_out;
SharedReg408_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg408_out;
SharedReg782_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg782_out;
SharedReg742_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg742_out;
SharedReg835_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg835_out;
SharedReg420_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg420_out;
SharedReg251_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg251_out;
SharedReg991_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg991_out;
   MUX_Product312_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg835_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg424_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg420_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg251_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg991_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg17_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay1No333_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg936_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg790_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg408_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg782_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg742_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg835_out_to_MUX_Product312_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product312_1_impl_0_out);

   Delay1No262_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product312_1_impl_0_out,
                 Y => Delay1No262_out);

SharedReg1284_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1284_out;
SharedReg1305_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1305_out;
SharedReg192_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg192_out;
SharedReg1263_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1263_out;
SharedReg993_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg993_out;
SharedReg1301_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1301_out;
SharedReg252_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg252_out;
SharedReg1278_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1278_out;
SharedReg1279_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1279_out;
SharedReg1292_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1292_out;
SharedReg1281_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1281_out;
SharedReg188_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg188_out;
SharedReg1059_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1059_out;
   MUX_Product312_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1284_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1305_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1281_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg188_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1059_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg192_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1263_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg993_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1301_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg252_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1278_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1279_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1292_out_to_MUX_Product312_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product312_1_impl_1_out);

   Delay1No263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product312_1_impl_1_out,
                 Y => Delay1No263_out);

Delay1No264_out_to_Product312_2_impl_parent_implementedSystem_port_0_cast <= Delay1No264_out;
Delay1No265_out_to_Product312_2_impl_parent_implementedSystem_port_1_cast <= Delay1No265_out;
   Product312_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product312_2_impl_out,
                 X => Delay1No264_out_to_Product312_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No265_out_to_Product312_2_impl_parent_implementedSystem_port_1_cast);

SharedReg427_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg427_out;
SharedReg851_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg851_out;
SharedReg843_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg843_out;
SharedReg1162_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1162_out;
SharedReg94_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg94_out;
SharedReg380_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg380_out;
SharedReg946_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg946_out;
SharedReg798_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg798_out;
SharedReg550_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg550_out;
SharedReg893_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg893_out;
SharedReg848_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg848_out;
SharedReg843_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg843_out;
SharedReg427_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg427_out;
   MUX_Product312_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg427_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg851_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg848_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg843_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg427_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg843_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1162_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg94_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg380_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg946_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg798_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg550_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg893_out_to_MUX_Product312_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product312_2_impl_0_out);

   Delay1No264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product312_2_impl_0_out,
                 Y => Delay1No264_out);

SharedReg1294_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1294_out;
SharedReg1311_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1311_out;
SharedReg1284_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1284_out;
SharedReg1285_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1285_out;
SharedReg269_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg269_out;
SharedReg1275_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1275_out;
SharedReg1005_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1005_out;
SharedReg1301_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1301_out;
SharedReg262_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg262_out;
SharedReg1278_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1278_out;
SharedReg1279_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1279_out;
SharedReg1292_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1292_out;
SharedReg1281_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1281_out;
   MUX_Product312_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1294_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1311_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1279_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1292_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1281_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1284_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1285_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg269_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1275_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1005_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1301_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg262_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1278_out_to_MUX_Product312_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product312_2_impl_1_out);

   Delay1No265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product312_2_impl_1_out,
                 Y => Delay1No265_out);

Delay1No266_out_to_Product312_3_impl_parent_implementedSystem_port_0_cast <= Delay1No266_out;
Delay1No267_out_to_Product312_3_impl_parent_implementedSystem_port_1_cast <= Delay1No267_out;
   Product312_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product312_3_impl_out,
                 X => Delay1No266_out_to_Product312_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No267_out_to_Product312_3_impl_parent_implementedSystem_port_1_cast);

SharedReg760_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg760_out;
SharedReg98_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg98_out;
SharedReg435_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg435_out;
SharedReg1171_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1171_out;
SharedReg905_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg905_out;
SharedReg102_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg102_out;
SharedReg104_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg104_out;
SharedReg387_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg387_out;
SharedReg1131_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1131_out;
SharedReg806_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg806_out;
SharedReg557_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg557_out;
SharedReg901_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg901_out;
SharedReg859_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg859_out;
   MUX_Product312_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg760_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg98_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg557_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg901_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg859_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg435_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1171_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg905_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg102_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg104_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg387_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1131_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg806_out_to_MUX_Product312_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product312_3_impl_0_out);

   Delay1No266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product312_3_impl_0_out,
                 Y => Delay1No266_out);

SharedReg1303_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1303_out;
SharedReg152_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg152_out;
SharedReg1294_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1294_out;
SharedReg1283_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1283_out;
SharedReg40_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg40_out;
SharedReg1040_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1040_out;
SharedReg279_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg279_out;
SharedReg1275_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1275_out;
SharedReg1096_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1096_out;
SharedReg1301_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1301_out;
SharedReg272_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg272_out;
SharedReg1278_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1278_out;
SharedReg1279_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1279_out;
   MUX_Product312_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1303_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg152_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg272_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1278_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1279_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1294_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1283_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg40_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1040_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg279_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1275_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1096_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1301_out_to_MUX_Product312_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product312_3_impl_1_out);

   Delay1No267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product312_3_impl_1_out,
                 Y => Delay1No267_out);

Delay1No268_out_to_Product312_4_impl_parent_implementedSystem_port_0_cast <= Delay1No268_out;
Delay1No269_out_to_Product312_4_impl_parent_implementedSystem_port_1_cast <= Delay1No269_out;
   Product312_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product312_4_impl_out,
                 X => Delay1No268_out_to_Product312_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No269_out_to_Product312_4_impl_parent_implementedSystem_port_1_cast);

SharedReg443_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg443_out;
SharedReg489_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg489_out;
SharedReg815_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg815_out;
SharedReg1076_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1076_out;
SharedReg767_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg767_out;
SharedReg1070_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1070_out;
SharedReg912_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg912_out;
SharedReg112_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg112_out;
SharedReg114_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg114_out;
SharedReg488_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg488_out;
SharedReg1073_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1073_out;
SharedReg868_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg868_out;
SharedReg566_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg566_out;
   MUX_Product312_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg443_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg489_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1073_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg868_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg566_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg815_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1076_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg767_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1070_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg912_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg112_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg114_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg488_out_to_MUX_Product312_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product312_4_impl_0_out);

   Delay1No268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product312_4_impl_0_out,
                 Y => Delay1No268_out);

SharedReg1290_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1290_out;
SharedReg1279_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1279_out;
SharedReg1303_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1303_out;
SharedReg343_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg343_out;
SharedReg1282_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1282_out;
SharedReg222_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg222_out;
SharedReg51_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg51_out;
SharedReg1124_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1124_out;
SharedReg289_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg289_out;
SharedReg1275_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1275_out;
SharedReg970_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg970_out;
SharedReg1301_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1301_out;
SharedReg282_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg282_out;
   MUX_Product312_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1290_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1279_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg970_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1301_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg282_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1303_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg343_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1282_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg222_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg51_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1124_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg289_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1275_out_to_MUX_Product312_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product312_4_impl_1_out);

   Delay1No269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product312_4_impl_1_out,
                 Y => Delay1No269_out);

Delay1No270_out_to_Product312_5_impl_parent_implementedSystem_port_0_cast <= Delay1No270_out;
Delay1No271_out_to_Product312_5_impl_parent_implementedSystem_port_1_cast <= Delay1No271_out;
   Product312_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product312_5_impl_out,
                 X => Delay1No270_out_to_Product312_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No271_out_to_Product312_5_impl_parent_implementedSystem_port_1_cast);

SharedReg346_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg346_out;
SharedReg1186_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1186_out;
SharedReg524_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg524_out;
SharedReg1208_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1208_out;
SharedReg916_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg916_out;
SharedReg821_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg821_out;
SharedReg1051_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1051_out;
SharedReg58_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg58_out;
SharedReg919_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg919_out;
SharedReg822_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg822_out;
SharedReg1259_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1259_out;
SharedReg63_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg63_out;
SharedReg55_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg55_out;
   MUX_Product312_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg346_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1186_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1259_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg63_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg55_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg524_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1208_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg916_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg821_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1051_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg58_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg919_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg822_out_to_MUX_Product312_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product312_5_impl_0_out);

   Delay1No270_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product312_5_impl_0_out,
                 Y => Delay1No270_out);

SharedReg167_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg167_out;
SharedReg1288_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1288_out;
SharedReg292_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg292_out;
SharedReg1290_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1290_out;
SharedReg1296_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1296_out;
SharedReg1309_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1309_out;
SharedReg1110_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1110_out;
SharedReg169_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg169_out;
SharedReg1283_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1283_out;
SharedReg1284_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1284_out;
SharedReg1285_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1285_out;
SharedReg295_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg295_out;
SharedReg166_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg166_out;
   MUX_Product312_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg167_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1288_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1285_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg295_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg166_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg292_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1290_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1296_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1309_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1110_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg169_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1283_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1284_out_to_MUX_Product312_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product312_5_impl_1_out);

   Delay1No271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product312_5_impl_1_out,
                 Y => Delay1No271_out);

Delay1No272_out_to_Product54_4_impl_parent_implementedSystem_port_0_cast <= Delay1No272_out;
Delay1No273_out_to_Product54_4_impl_parent_implementedSystem_port_1_cast <= Delay1No273_out;
   Product54_4_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product54_4_impl_out,
                 X => Delay1No272_out_to_Product54_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No273_out_to_Product54_4_impl_parent_implementedSystem_port_1_cast);

SharedReg907_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg907_out;
SharedReg867_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg867_out;
SharedReg862_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg862_out;
SharedReg108_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg108_out;
SharedReg47_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg47_out;
SharedReg1179_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1179_out;
SharedReg910_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg910_out;
SharedReg975_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg975_out;
SharedReg52_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg52_out;
SharedReg44_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg44_out;
SharedReg337_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_11_cast <= SharedReg337_out;
Delay20No16_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_12_cast <= Delay20No16_out;
SharedReg610_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg610_out;
   MUX_Product54_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg907_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg867_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg337_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay20No16_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg610_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg862_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg108_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg47_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1179_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg910_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg975_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg52_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg44_out_to_MUX_Product54_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product54_4_impl_0_out);

   Delay1No272_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product54_4_impl_0_out,
                 Y => Delay1No272_out);

SharedReg1278_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1278_out;
SharedReg1279_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1279_out;
SharedReg1292_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1292_out;
SharedReg160_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg160_out;
SharedReg161_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_5_cast <= SharedReg161_out;
SharedReg1283_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1283_out;
SharedReg1284_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1284_out;
SharedReg165_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg165_out;
SharedReg285_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg285_out;
SharedReg158_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg158_out;
SharedReg159_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg159_out;
SharedReg1297_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1297_out;
SharedReg163_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg163_out;
   MUX_Product54_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1278_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1279_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg159_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1297_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg163_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1292_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg160_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg161_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1283_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1284_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg165_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg285_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg158_out_to_MUX_Product54_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product54_4_impl_1_out);

   Delay1No273_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product54_4_impl_1_out,
                 Y => Delay1No273_out);

Delay1No274_out_to_Product54_5_impl_parent_implementedSystem_port_0_cast <= Delay1No274_out;
Delay1No275_out_to_Product54_5_impl_parent_implementedSystem_port_1_cast <= Delay1No275_out;
   Product54_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product54_5_impl_out,
                 X => Delay1No274_out_to_Product54_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No275_out_to_Product54_5_impl_parent_implementedSystem_port_1_cast);

SharedReg1189_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1189_out;
SharedReg1201_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1201_out;
SharedReg573_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg573_out;
SharedReg871_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg871_out;
SharedReg1204_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1204_out;
SharedReg1203_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1203_out;
SharedReg1051_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1051_out;
SharedReg293_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg293_out;
SharedReg917_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg917_out;
SharedReg120_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg120_out;
SharedReg1262_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1262_out;
SharedReg1186_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg1186_out;
Delay1No337_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_13_cast <= Delay1No337_out;
   MUX_Product54_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1189_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1201_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1262_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1186_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => Delay1No337_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg573_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg871_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1204_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1203_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1051_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg293_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg917_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg120_out_to_MUX_Product54_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product54_5_impl_0_out);

   Delay1No274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product54_5_impl_0_out,
                 Y => Delay1No274_out);

SharedReg1276_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1276_out;
SharedReg1288_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1288_out;
SharedReg171_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg171_out;
SharedReg1278_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1278_out;
SharedReg1291_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1291_out;
SharedReg1280_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1280_out;
SharedReg352_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg352_out;
SharedReg1111_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1111_out;
SharedReg1283_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1283_out;
SharedReg1105_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1105_out;
SharedReg1305_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1305_out;
SharedReg1295_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1295_out;
SharedReg1263_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1263_out;
   MUX_Product54_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1276_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1288_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1305_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1295_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1263_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg171_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1278_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1291_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1280_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg352_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1111_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1283_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1105_out_to_MUX_Product54_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Product54_5_impl_1_out);

   Delay1No275_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product54_5_impl_1_out,
                 Y => Delay1No275_out);

Delay1No276_out_to_Product62_5_impl_parent_implementedSystem_port_0_cast <= Delay1No276_out;
Delay1No277_out_to_Product62_5_impl_parent_implementedSystem_port_1_cast <= Delay1No277_out;
   Product62_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product62_5_impl_out,
                 X => Delay1No276_out_to_Product62_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No277_out_to_Product62_5_impl_parent_implementedSystem_port_1_cast);

SharedReg61_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg61_out;
SharedReg59_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg59_out;
SharedReg118_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg118_out;
Delay1No343_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_4_cast <= Delay1No343_out;
SharedReg769_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg769_out;
SharedReg1184_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1184_out;
SharedReg1200_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1200_out;
SharedReg920_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg920_out;
Delay64No5_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_9_cast <= Delay64No5_out;
SharedReg1208_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1208_out;
SharedReg1259_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg1259_out;
SharedReg913_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg913_out;
   MUX_Product62_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg61_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg59_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1259_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg913_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg118_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => Delay1No343_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg769_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1184_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1200_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg920_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => Delay64No5_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1208_out_to_MUX_Product62_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product62_5_impl_0_LUT_out,
                 oMux => MUX_Product62_5_impl_0_out);

   Delay1No276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product62_5_impl_0_out,
                 Y => Delay1No276_out);

SharedReg65_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg65_out;
SharedReg168_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg168_out;
SharedReg236_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg236_out;
SharedReg1249_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1249_out;
SharedReg1279_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1279_out;
SharedReg1314_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1314_out;
SharedReg1278_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1278_out;
SharedReg1311_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1311_out;
SharedReg1294_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1294_out;
SharedReg1284_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1284_out;
SharedReg1303_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1303_out;
SharedReg1263_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1263_out;
   MUX_Product62_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_12_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg65_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg168_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1303_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1263_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_2 => SharedReg236_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1249_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1279_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1314_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1278_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1311_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1294_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1284_out_to_MUX_Product62_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product62_5_impl_1_LUT_out,
                 oMux => MUX_Product62_5_impl_1_out);

   Delay1No277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product62_5_impl_1_out,
                 Y => Delay1No277_out);

Delay1No278_out_to_Subtract12_0_impl_parent_implementedSystem_port_0_cast <= Delay1No278_out;
Delay1No279_out_to_Subtract12_0_impl_parent_implementedSystem_port_1_cast <= Delay1No279_out;
   Subtract12_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_0_impl_out,
                 X => Delay1No278_out_to_Subtract12_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No279_out_to_Subtract12_0_impl_parent_implementedSystem_port_1_cast);

SharedReg587_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg587_out;
SharedReg454_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg454_out;
Delay84No_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_3_cast <= Delay84No_out;
SharedReg360_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg360_out;
SharedReg534_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg534_out;
SharedReg680_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg680_out;
SharedReg780_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg780_out;
SharedReg362_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg362_out;
SharedReg533_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg533_out;
SharedReg676_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg676_out;
Delay48No_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_11_cast <= Delay48No_out;
SharedReg401_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg401_out;
SharedReg628_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg628_out;
   MUX_Subtract12_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg587_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg454_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay48No_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg401_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg628_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => Delay84No_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg360_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg534_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg680_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg780_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg362_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg533_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg676_out_to_MUX_Subtract12_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract12_0_impl_0_out);

   Delay1No278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_0_impl_0_out,
                 Y => Delay1No278_out);

Delay73No_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_1_cast <= Delay73No_out;
SharedReg1086_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1086_out;
SharedReg1084_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1084_out;
SharedReg1147_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1147_out;
SharedReg977_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg977_out;
SharedReg931_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg931_out;
SharedReg928_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg928_out;
SharedReg924_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg924_out;
SharedReg924_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg924_out;
SharedReg1140_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1140_out;
SharedReg924_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg924_out;
SharedReg980_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg980_out;
SharedReg924_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg924_out;
   MUX_Subtract12_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay73No_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1086_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg924_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg980_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg924_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1084_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1147_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg977_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg931_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg928_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg924_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg924_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1140_out_to_MUX_Subtract12_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract12_0_impl_1_out);

   Delay1No279_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_0_impl_1_out,
                 Y => Delay1No279_out);

Delay1No280_out_to_Subtract12_1_impl_parent_implementedSystem_port_0_cast <= Delay1No280_out;
Delay1No281_out_to_Subtract12_1_impl_parent_implementedSystem_port_1_cast <= Delay1No281_out;
   Subtract12_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_1_impl_out,
                 X => Delay1No280_out_to_Subtract12_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No281_out_to_Subtract12_1_impl_parent_implementedSystem_port_1_cast);

SharedReg409_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg409_out;
SharedReg635_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg635_out;
SharedReg688_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg688_out;
SharedReg460_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg460_out;
Delay84No1_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_5_cast <= Delay84No1_out;
SharedReg367_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg367_out;
SharedReg543_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg543_out;
SharedReg687_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg687_out;
SharedReg788_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg788_out;
SharedReg370_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg370_out;
SharedReg685_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg685_out;
SharedReg684_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg684_out;
SharedReg377_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg377_out;
   MUX_Subtract12_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg409_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg635_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg685_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg684_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg377_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg688_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg460_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay84No1_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg367_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg543_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg687_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg788_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg370_out_to_MUX_Subtract12_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract12_1_impl_0_out);

   Delay1No280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_1_impl_0_out,
                 Y => Delay1No280_out);

SharedReg994_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg994_out;
SharedReg977_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg977_out;
SharedReg989_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg989_out;
SharedReg1062_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1062_out;
SharedReg935_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg935_out;
Delay79No1_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_6_cast <= Delay79No1_out;
SharedReg991_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg991_out;
SharedReg988_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg988_out;
SharedReg983_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg983_out;
SharedReg933_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg933_out;
SharedReg933_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg933_out;
SharedReg1061_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1061_out;
SharedReg977_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg977_out;
   MUX_Subtract12_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg994_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg977_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg933_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1061_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg977_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg989_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1062_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg935_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => Delay79No1_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg991_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg988_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg983_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg933_out_to_MUX_Subtract12_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract12_1_impl_1_out);

   Delay1No281_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_1_impl_1_out,
                 Y => Delay1No281_out);

Delay1No282_out_to_Subtract12_2_impl_parent_implementedSystem_port_0_cast <= Delay1No282_out;
Delay1No283_out_to_Subtract12_2_impl_parent_implementedSystem_port_1_cast <= Delay1No283_out;
   Subtract12_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_2_impl_out,
                 X => Delay1No282_out_to_Subtract12_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No283_out_to_Subtract12_2_impl_parent_implementedSystem_port_1_cast);

SharedReg690_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg690_out;
Delay48No2_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_2_cast <= Delay48No2_out;
SharedReg419_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg419_out;
SharedReg643_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg643_out;
SharedReg695_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg695_out;
SharedReg510_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg510_out;
Delay84No2_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_7_cast <= Delay84No2_out;
SharedReg374_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg374_out;
SharedReg601_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg601_out;
SharedReg751_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg751_out;
SharedReg795_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg795_out;
SharedReg378_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg378_out;
SharedReg691_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg691_out;
   MUX_Subtract12_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg690_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay48No2_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg795_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg378_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg691_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg419_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg643_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg695_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg510_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => Delay84No2_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg374_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg601_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg751_out_to_MUX_Subtract12_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract12_2_impl_0_out);

   Delay1No282_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_2_impl_0_out,
                 Y => Delay1No282_out);

SharedReg1004_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1004_out;
SharedReg991_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg991_out;
SharedReg959_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg959_out;
SharedReg1017_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1017_out;
SharedReg953_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg953_out;
SharedReg1021_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1021_out;
SharedReg1092_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1092_out;
Delay79No2_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_8_cast <= Delay79No2_out;
SharedReg1002_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1002_out;
SharedReg962_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg962_out;
SharedReg950_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg950_out;
SharedReg943_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg943_out;
SharedReg943_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg943_out;
   MUX_Subtract12_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1004_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg991_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg950_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg943_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg943_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg959_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1017_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg953_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1021_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1092_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => Delay79No2_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1002_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg962_out_to_MUX_Subtract12_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract12_2_impl_1_out);

   Delay1No283_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_2_impl_1_out,
                 Y => Delay1No283_out);

Delay1No284_out_to_Subtract12_3_impl_parent_implementedSystem_port_0_cast <= Delay1No284_out;
Delay1No285_out_to_Subtract12_3_impl_parent_implementedSystem_port_1_cast <= Delay1No285_out;
   Subtract12_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_3_impl_out,
                 X => Delay1No284_out_to_Subtract12_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No285_out_to_Subtract12_3_impl_parent_implementedSystem_port_1_cast);

SharedReg432_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg432_out;
SharedReg702_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg702_out;
SharedReg700_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg700_out;
SharedReg522_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg522_out;
SharedReg426_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg426_out;
SharedReg701_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg701_out;
SharedReg705_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg705_out;
SharedReg515_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg515_out;
SharedReg565_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg565_out;
SharedReg382_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg382_out;
SharedReg609_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg609_out;
SharedReg759_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg759_out;
SharedReg857_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg857_out;
   MUX_Subtract12_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg432_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg702_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg609_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg759_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg857_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg700_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg522_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg426_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg701_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg705_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg515_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg565_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg382_out_to_MUX_Subtract12_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract12_3_impl_0_out);

   Delay1No284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_3_impl_0_out,
                 Y => Delay1No284_out);

SharedReg956_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg956_out;
SharedReg956_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg956_out;
SharedReg1130_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1130_out;
SharedReg1091_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1091_out;
SharedReg1032_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1032_out;
SharedReg1028_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1028_out;
SharedReg964_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg964_out;
SharedReg1093_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1093_out;
SharedReg1095_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1095_out;
SharedReg1102_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1102_out;
SharedReg1028_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1028_out;
SharedReg1038_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1038_out;
SharedReg960_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg960_out;
   MUX_Subtract12_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg956_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg956_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1028_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1038_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg960_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1130_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1091_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1032_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1028_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg964_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1093_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1095_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1102_out_to_MUX_Subtract12_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract12_3_impl_1_out);

   Delay1No285_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_3_impl_1_out,
                 Y => Delay1No285_out);

Delay1No286_out_to_Subtract12_4_impl_parent_implementedSystem_port_0_cast <= Delay1No286_out;
Delay1No287_out_to_Subtract12_4_impl_parent_implementedSystem_port_1_cast <= Delay1No287_out;
   Subtract12_4_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_4_impl_out,
                 X => Delay1No286_out_to_Subtract12_4_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No287_out_to_Subtract12_4_impl_parent_implementedSystem_port_1_cast);

SharedReg911_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_1_cast <= SharedReg911_out;
SharedReg866_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_2_cast <= SharedReg866_out;
SharedReg486_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_3_cast <= SharedReg486_out;
SharedReg711_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_4_cast <= SharedReg711_out;
SharedReg762_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_5_cast <= SharedReg762_out;
SharedReg492_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_6_cast <= SharedReg492_out;
SharedReg480_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_7_cast <= SharedReg480_out;
SharedReg710_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_8_cast <= SharedReg710_out;
SharedReg713_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_9_cast <= SharedReg713_out;
SharedReg668_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_10_cast <= SharedReg668_out;
Delay84No4_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_11_cast <= Delay84No4_out;
SharedReg439_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_12_cast <= SharedReg439_out;
SharedReg765_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_13_cast <= SharedReg765_out;
   MUX_Subtract12_4_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg911_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg866_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => Delay84No4_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg439_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg765_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg486_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg711_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg762_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg492_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg480_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg710_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg713_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg668_out_to_MUX_Subtract12_4_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract12_4_impl_0_out);

   Delay1No286_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_4_impl_0_out,
                 Y => Delay1No286_out);

Delay58No4_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_1_cast <= Delay58No4_out;
SharedReg1035_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1035_out;
SharedReg1028_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1028_out;
SharedReg965_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_4_cast <= SharedReg965_out;
Delay5No22_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_5_cast <= Delay5No22_out;
SharedReg1011_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1011_out;
SharedReg1013_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1013_out;
SharedReg1011_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1011_out;
SharedReg1042_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1042_out;
SharedReg1013_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1013_out;
SharedReg1072_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1072_out;
Delay79No4_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_12_cast <= Delay79No4_out;
SharedReg1011_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1011_out;
   MUX_Subtract12_4_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay58No4_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1035_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1072_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => Delay79No4_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1011_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg1028_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg965_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => Delay5No22_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1011_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1013_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1011_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1042_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1013_out_to_MUX_Subtract12_4_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract12_4_impl_1_out);

   Delay1No287_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_4_impl_1_out,
                 Y => Delay1No287_out);

Delay1No288_out_to_Subtract12_5_impl_parent_implementedSystem_port_0_cast <= Delay1No288_out;
Delay1No289_out_to_Subtract12_5_impl_parent_implementedSystem_port_1_cast <= Delay1No289_out;
   Subtract12_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_true_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Subtract12_5_impl_out,
                 X => Delay1No288_out_to_Subtract12_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No289_out_to_Subtract12_5_impl_parent_implementedSystem_port_1_cast);

Delay84No5_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_1_cast <= Delay84No5_out;
SharedReg444_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_2_cast <= SharedReg444_out;
SharedReg721_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg721_out;
SharedReg876_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg876_out;
SharedReg1188_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1188_out;
SharedReg530_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg530_out;
SharedReg671_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg671_out;
SharedReg769_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg769_out;
SharedReg1261_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1261_out;
SharedReg574_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg574_out;
SharedReg820_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_11_cast <= SharedReg820_out;
SharedReg622_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_12_cast <= SharedReg622_out;
SharedReg624_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_13_cast <= SharedReg624_out;
   MUX_Subtract12_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay84No5_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg444_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg820_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg622_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg624_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg721_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg876_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1188_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg530_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg671_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg769_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1261_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg574_out_to_MUX_Subtract12_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract12_5_impl_0_out);

   Delay1No288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_5_impl_0_out,
                 Y => Delay1No288_out);

SharedReg1106_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1106_out;
SharedReg1126_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1126_out;
SharedReg968_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg968_out;
SharedReg1055_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1055_out;
SharedReg1122_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1122_out;
SharedReg1044_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1044_out;
SharedReg968_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg968_out;
SharedReg1047_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1047_out;
SharedReg968_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg968_out;
SharedReg1108_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1108_out;
SharedReg1044_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_11_cast <= SharedReg1044_out;
SharedReg1057_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_12_cast <= SharedReg1057_out;
SharedReg1049_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_13_cast <= SharedReg1049_out;
   MUX_Subtract12_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_13_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1106_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1126_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg1044_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg1057_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg1049_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_13_cast,
                 iS_2 => SharedReg968_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1055_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1122_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1044_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg968_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1047_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg968_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1108_out_to_MUX_Subtract12_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount131_out,
                 oMux => MUX_Subtract12_5_impl_1_out);

   Delay1No289_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Subtract12_5_impl_1_out,
                 Y => Delay1No289_out);

Delay1No290_out_to_Add10_5_impl_parent_implementedSystem_port_0_cast <= Delay1No290_out;
Delay1No291_out_to_Add10_5_impl_parent_implementedSystem_port_1_cast <= Delay1No291_out;
   Add10_5_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Add10_5_impl_out,
                 X => Delay1No290_out_to_Add10_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No291_out_to_Add10_5_impl_parent_implementedSystem_port_1_cast);

Delay5No17_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_1_cast <= Delay5No17_out;
Delay60No5_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_2_cast <= Delay60No5_out;
Delay55No11_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_3_cast <= Delay55No11_out;
SharedReg1208_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1208_out;
SharedReg871_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg871_out;
SharedReg918_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg918_out;
SharedReg1206_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1206_out;
SharedReg1202_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg1202_out;
SharedReg1185_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1185_out;
SharedReg1205_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1205_out;
   MUX_Add10_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_10_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => Delay5No17_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay60No5_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay55No11_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1208_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg871_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg918_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1206_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1202_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1185_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1205_out_to_MUX_Add10_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add10_5_impl_0_LUT_out,
                 oMux => MUX_Add10_5_impl_0_out);

   Delay1No290_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add10_5_impl_0_out,
                 Y => Delay1No290_out);

SharedReg1104_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg1104_out;
SharedReg1248_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1248_out;
SharedReg1248_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1248_out;
SharedReg1248_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1248_out;
SharedReg1104_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1104_out;
SharedReg1248_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1248_out;
SharedReg1248_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1248_out;
SharedReg1248_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1248_out;
SharedReg1242_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1242_out;
SharedReg1257_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1257_out;
   MUX_Add10_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_10_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1104_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1248_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1248_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1248_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1104_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1248_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1248_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1248_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1242_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1257_out_to_MUX_Add10_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Add10_5_impl_1_LUT_out,
                 oMux => MUX_Add10_5_impl_1_out);

   Delay1No291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Add10_5_impl_1_out,
                 Y => Delay1No291_out);
   Constant1_0_impl_instance: Constant_float_8_23_1_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_0_impl_out);

Delay1No292_out_to_Divide_0_impl_parent_implementedSystem_port_0_cast <= Delay1No292_out;
Delay1No293_out_to_Divide_0_impl_parent_implementedSystem_port_1_cast <= Delay1No293_out;
   Divide_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_div_Y_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Divide_0_impl_out,
                 X => Delay1No292_out_to_Divide_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No293_out_to_Divide_0_impl_parent_implementedSystem_port_1_cast);

SharedReg1255_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg1255_out;
SharedReg1255_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg1255_out;
SharedReg1255_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg1255_out;
SharedReg1255_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1255_out;
SharedReg1255_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1255_out;
SharedReg1255_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg1255_out;
   MUX_Divide_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg1255_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1255_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1255_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1255_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1255_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1255_out_to_MUX_Divide_0_impl_0_parent_implementedSystem_port_6_cast,
                 iSel => MUX_Divide_0_impl_0_LUT_out,
                 oMux => MUX_Divide_0_impl_0_out);

   Delay1No292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Divide_0_impl_0_out,
                 Y => Delay1No292_out);

SharedReg977_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg977_out;
SharedReg1017_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1017_out;
SharedReg1091_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1091_out;
SharedReg965_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg965_out;
SharedReg1115_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1115_out;
SharedReg968_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg968_out;
   MUX_Divide_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_6_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg977_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1017_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1091_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg965_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1115_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg968_out_to_MUX_Divide_0_impl_1_parent_implementedSystem_port_6_cast,
                 iSel => MUX_Divide_0_impl_1_LUT_out,
                 oMux => MUX_Divide_0_impl_1_out);

   Delay1No293_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Divide_0_impl_1_out,
                 Y => Delay1No293_out);

Delay1No294_out_to_Product213_5_impl_parent_implementedSystem_port_0_cast <= Delay1No294_out;
Delay1No295_out_to_Product213_5_impl_parent_implementedSystem_port_1_cast <= Delay1No295_out;
   Product213_5_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product213_5_impl_out,
                 X => Delay1No294_out_to_Product213_5_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No295_out_to_Product213_5_impl_parent_implementedSystem_port_1_cast);

SharedReg291_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_1_cast <= SharedReg291_out;
Delay1No349_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_2_cast <= Delay1No349_out;
SharedReg915_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_3_cast <= SharedReg915_out;
SharedReg1185_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_4_cast <= SharedReg1185_out;
SharedReg1201_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_5_cast <= SharedReg1201_out;
SharedReg769_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_6_cast <= SharedReg769_out;
SharedReg1208_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_7_cast <= SharedReg1208_out;
SharedReg824_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_8_cast <= SharedReg824_out;
SharedReg1183_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_9_cast <= SharedReg1183_out;
SharedReg1248_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_10_cast <= SharedReg1248_out;
   MUX_Product213_5_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_10_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg291_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay1No349_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg915_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1185_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1201_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg769_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1208_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg824_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1183_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1248_out_to_MUX_Product213_5_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product213_5_impl_0_LUT_out,
                 oMux => MUX_Product213_5_impl_0_out);

   Delay1No294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_5_impl_0_out,
                 Y => Delay1No294_out);

SharedReg232_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_1_cast <= SharedReg232_out;
SharedReg1104_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_2_cast <= SharedReg1104_out;
SharedReg1274_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_3_cast <= SharedReg1274_out;
SharedReg1279_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_4_cast <= SharedReg1279_out;
SharedReg1281_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_5_cast <= SharedReg1281_out;
SharedReg1266_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_6_cast <= SharedReg1266_out;
SharedReg1292_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_7_cast <= SharedReg1292_out;
SharedReg1272_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_8_cast <= SharedReg1272_out;
SharedReg1289_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_9_cast <= SharedReg1289_out;
SharedReg1263_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_10_cast <= SharedReg1263_out;
   MUX_Product213_5_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_10_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg232_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg1104_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg1274_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg1279_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg1281_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg1266_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg1292_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg1272_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg1289_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg1263_out_to_MUX_Product213_5_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product213_5_impl_1_LUT_out,
                 oMux => MUX_Product213_5_impl_1_out);

   Delay1No295_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product213_5_impl_1_out,
                 Y => Delay1No295_out);
   Constant_0_impl_instance: Constant_float_8_23_348_mult_8en9_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_0_impl_out);

   Delay5No_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UU_del_1_0_out,
                 Y => Delay5No_out);

   Delay5No1_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UU_del_1_1_out,
                 Y => Delay5No1_out);

   Delay5No2_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UU_del_1_2_out,
                 Y => Delay5No2_out);

   Delay5No3_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UU_del_1_3_out,
                 Y => Delay5No3_out);

   Delay5No4_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UU_del_1_4_out,
                 Y => Delay5No4_out);

   Delay5No5_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UU_del_1_5_out,
                 Y => Delay5No5_out);

   Delay90No_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg10_out,
                 Y => Delay90No_out);

   Delay90No1_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg21_out,
                 Y => Delay90No1_out);

   Delay90No2_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => Delay90No2_out);

   Delay90No3_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => Delay90No3_out);

   Delay90No4_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => Delay90No4_out);

   Delay90No5_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => Delay90No5_out);

   Delay102No_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => Delay102No_out);

   Delay102No1_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg85_out,
                 Y => Delay102No1_out);

   Delay102No2_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg95_out,
                 Y => Delay102No2_out);

   Delay102No3_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg105_out,
                 Y => Delay102No3_out);

   Delay102No4_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg115_out,
                 Y => Delay102No4_out);

   Delay102No5_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg125_out,
                 Y => Delay102No5_out);

   Delay94No_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => Delay94No_out);

   Delay94No1_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg141_out,
                 Y => Delay94No1_out);

   Delay94No2_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => Delay94No2_out);

   Delay94No3_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg157_out,
                 Y => Delay94No3_out);

   Delay94No4_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => Delay94No4_out);

   Delay94No5_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg173_out,
                 Y => Delay94No5_out);

   Delay5No6_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VV_del_1_0_out,
                 Y => Delay5No6_out);

   Delay5No7_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VV_del_1_1_out,
                 Y => Delay5No7_out);

   Delay5No8_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VV_del_1_2_out,
                 Y => Delay5No8_out);

   Delay5No9_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VV_del_1_3_out,
                 Y => Delay5No9_out);

   Delay5No10_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VV_del_1_4_out,
                 Y => Delay5No10_out);

   Delay5No11_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VV_del_1_5_out,
                 Y => Delay5No11_out);

   Delay102No6_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg184_out,
                 Y => Delay102No6_out);

   Delay102No7_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg195_out,
                 Y => Delay102No7_out);

   Delay102No8_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg206_out,
                 Y => Delay102No8_out);

   Delay102No9_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg217_out,
                 Y => Delay102No9_out);

   Delay102No10_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg228_out,
                 Y => Delay102No10_out);

   Delay102No11_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg239_out,
                 Y => Delay102No11_out);

   Delay97No_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg249_out,
                 Y => Delay97No_out);

   Delay97No1_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg259_out,
                 Y => Delay97No1_out);

   Delay97No2_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg269_out,
                 Y => Delay97No2_out);

   Delay97No3_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg279_out,
                 Y => Delay97No3_out);

   Delay97No4_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg289_out,
                 Y => Delay97No4_out);

   Delay97No5_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg299_out,
                 Y => Delay97No5_out);

   Delay78No6_instance: Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=50 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg308_out,
                 Y => Delay78No6_out);

   Delay78No7_instance: Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=50 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg317_out,
                 Y => Delay78No7_out);

   Delay78No8_instance: Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=50 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg326_out,
                 Y => Delay78No8_out);

   Delay78No9_instance: Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=50 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg335_out,
                 Y => Delay78No9_out);

   Delay78No10_instance: Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=50 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg344_out,
                 Y => Delay78No10_out);

   Delay78No11_instance: Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=50 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg353_out,
                 Y => Delay78No11_out);

   Delay5No12_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WW_del_1_0_out,
                 Y => Delay5No12_out);

   Delay5No13_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WW_del_1_1_out,
                 Y => Delay5No13_out);

   Delay5No14_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WW_del_1_2_out,
                 Y => Delay5No14_out);

   Delay5No15_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WW_del_1_3_out,
                 Y => Delay5No15_out);

   Delay5No16_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WW_del_1_4_out,
                 Y => Delay5No16_out);

   Delay5No17_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WW_del_1_5_out,
                 Y => Delay5No17_out);

   Delay1No332_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_U_0_out,
                 Y => Delay1No332_out);

   Delay1No333_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_U_1_out,
                 Y => Delay1No333_out);

   Delay1No334_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_U_2_out,
                 Y => Delay1No334_out);

   Delay1No335_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_U_3_out,
                 Y => Delay1No335_out);

   Delay1No336_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_U_4_out,
                 Y => Delay1No336_out);

   Delay1No337_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_U_5_out,
                 Y => Delay1No337_out);

   Delay1No338_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_V_0_out,
                 Y => Delay1No338_out);

   Delay1No339_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_V_1_out,
                 Y => Delay1No339_out);

   Delay1No340_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_V_2_out,
                 Y => Delay1No340_out);

   Delay1No341_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_V_3_out,
                 Y => Delay1No341_out);

   Delay1No342_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_V_4_out,
                 Y => Delay1No342_out);

   Delay1No343_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_V_5_out,
                 Y => Delay1No343_out);

   Delay1No344_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_W_0_out,
                 Y => Delay1No344_out);

   Delay1No345_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_W_1_out,
                 Y => Delay1No345_out);

   Delay1No346_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_W_2_out,
                 Y => Delay1No346_out);

   Delay1No347_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_W_3_out,
                 Y => Delay1No347_out);

   Delay1No348_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_W_4_out,
                 Y => Delay1No348_out);

   Delay1No349_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => R_W_5_out,
                 Y => Delay1No349_out);

   Delay58No4_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1016_out,
                 Y => Delay58No4_out);

   Delay73No_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg932_out,
                 Y => Delay73No_out);

   Delay5No22_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg967_out,
                 Y => Delay5No22_out);

   Delay79No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg955_out,
                 Y => Delay79No1_out);

   Delay79No2_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg964_out,
                 Y => Delay79No2_out);

   Delay79No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1081_out,
                 Y => Delay79No4_out);

   Delay9No39_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1093_out,
                 Y => Delay9No39_out);

   Delay88No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg362_out,
                 Y => Delay88No_out);

   Delay88No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg370_out,
                 Y => Delay88No1_out);

   Delay88No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg378_out,
                 Y => Delay88No2_out);

   Delay88No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg432_out,
                 Y => Delay88No3_out);

   Delay88No4_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg441_out,
                 Y => Delay88No4_out);

   Delay88No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg530_out,
                 Y => Delay88No5_out);

   Delay76No3_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg516_out,
                 Y => Delay76No3_out);

   Delay6No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg609_out,
                 Y => Delay6No3_out);

   Delay87No8_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg470_out,
                 Y => Delay87No8_out);

   Delay87No9_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg565_out,
                 Y => Delay87No9_out);

   Delay87No10_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg572_out,
                 Y => Delay87No10_out);

   Delay87No11_instance: Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=39 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg492_out,
                 Y => Delay87No11_out);

   Delay96No_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg407_out,
                 Y => Delay96No_out);

   Delay96No1_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg417_out,
                 Y => Delay96No1_out);

   Delay96No2_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg424_out,
                 Y => Delay96No2_out);

   Delay96No3_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg478_out,
                 Y => Delay96No3_out);

   Delay96No4_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg486_out,
                 Y => Delay96No4_out);

   Delay96No5_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg580_out,
                 Y => Delay96No5_out);

   Delay62No_instance: Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=42 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg455_out,
                 Y => Delay62No_out);

   Delay104No_instance: Delay_34_DelayLength_95_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=95 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg588_out,
                 Y => Delay104No_out);

   Delay104No1_instance: Delay_34_DelayLength_87_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=87 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg596_out,
                 Y => Delay104No1_out);

   Delay104No2_instance: Delay_34_DelayLength_85_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=85 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg651_out,
                 Y => Delay104No2_out);

   Delay104No3_instance: Delay_34_DelayLength_85_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=85 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg660_out,
                 Y => Delay104No3_out);

   Delay104No5_instance: Delay_34_DelayLength_97_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=97 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg774_out,
                 Y => Delay104No5_out);

   Delay67No4_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg523_out,
                 Y => Delay67No4_out);

   Delay24No1_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg503_out,
                 Y => Delay24No1_out);

   Delay24No2_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg510_out,
                 Y => Delay24No2_out);

   Delay78No18_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg683_out,
                 Y => Delay78No18_out);

   Delay78No19_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg842_out,
                 Y => Delay78No19_out);

   Delay78No20_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg851_out,
                 Y => Delay78No20_out);

   Delay19No7_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg641_out,
                 Y => Delay19No7_out);

   Delay19No10_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg668_out,
                 Y => Delay19No10_out);

   Delay73No6_instance: Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=49 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg498_out,
                 Y => Delay73No6_out);

   Delay73No8_instance: Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=64 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg604_out,
                 Y => Delay73No8_out);

   Delay73No9_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg708_out,
                 Y => Delay73No9_out);

   Delay73No10_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg717_out,
                 Y => Delay73No10_out);

   Delay73No11_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg626_out,
                 Y => Delay73No11_out);

   Delay84No_instance: Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=65 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg539_out,
                 Y => Delay84No_out);

   Delay84No1_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg549_out,
                 Y => Delay84No1_out);

   Delay84No2_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg556_out,
                 Y => Delay84No2_out);

   Delay84No4_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg617_out,
                 Y => Delay84No4_out);

   Delay84No5_instance: Delay_34_DelayLength_68_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=68 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg725_out,
                 Y => Delay84No5_out);

   Delay14No4_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg399_out,
                 Y => Delay14No4_out);

   Delay104No6_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg734_out,
                 Y => Delay104No6_out);

   Delay104No7_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg745_out,
                 Y => Delay104No7_out);

   Delay104No8_instance: Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=45 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg754_out,
                 Y => Delay104No8_out);

   Delay104No9_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg808_out,
                 Y => Delay104No9_out);

   Delay104No11_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg923_out,
                 Y => Delay104No11_out);

   Delay88No6_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg633_out,
                 Y => Delay88No6_out);

   Delay88No7_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg689_out,
                 Y => Delay88No7_out);

   Delay88No8_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg699_out,
                 Y => Delay88No8_out);

   Delay88No9_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg861_out,
                 Y => Delay88No9_out);

   Delay88No10_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg870_out,
                 Y => Delay88No10_out);

   Delay88No11_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg826_out,
                 Y => Delay88No11_out);

   Delay59No5_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg675_out,
                 Y => Delay59No5_out);

   Delay76No7_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg790_out,
                 Y => Delay76No7_out);

   Delay76No9_instance: Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=57 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1173_out,
                 Y => Delay76No9_out);

   Delay89No8_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg799_out,
                 Y => Delay89No8_out);

   Delay89No10_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1182_out,
                 Y => Delay89No10_out);

   Delay69No10_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg768_out,
                 Y => Delay69No10_out);

   Delay69No11_instance: Delay_34_DelayLength_61_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=61 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg878_out,
                 Y => Delay69No11_out);

   Delay70No_instance: Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=64 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1217_out,
                 Y => Delay70No_out);

   Delay70No1_instance: Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=64 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1223_out,
                 Y => Delay70No1_out);

   Delay70No2_instance: Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=64 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1229_out,
                 Y => Delay70No2_out);

   Delay70No3_instance: Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=64 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1235_out,
                 Y => Delay70No3_out);

   Delay70No4_instance: Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=64 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1241_out,
                 Y => Delay70No4_out);

   Delay70No5_instance: Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=64 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1247_out,
                 Y => Delay70No5_out);

   Delay60No_instance: Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=40 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg781_out,
                 Y => Delay60No_out);

   Delay60No3_instance: Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=50 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg393_out,
                 Y => Delay60No3_out);

   Delay60No4_instance: Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=50 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1199_out,
                 Y => Delay60No4_out);

   Delay60No5_instance: Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=40 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1190_out,
                 Y => Delay60No5_out);

   Delay55No6_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg886_out,
                 Y => Delay55No6_out);

   Delay55No7_instance: Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=43 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1159_out,
                 Y => Delay55No7_out);

   Delay55No8_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1166_out,
                 Y => Delay55No8_out);

   Delay55No11_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1211_out,
                 Y => Delay55No11_out);

   Delay69No12_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg462_out,
                 Y => Delay69No12_out);

   Delay20No16_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg912_out,
                 Y => Delay20No16_out);

   Delay48No_instance: Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=42 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1152_out,
                 Y => Delay48No_out);

   Delay48No2_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg385_out,
                 Y => Delay48No2_out);

   Delay19No13_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg892_out,
                 Y => Delay19No13_out);

   Delay64No_instance: Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=44 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg834_out,
                 Y => Delay64No_out);

   Delay64No3_instance: Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=49 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg906_out,
                 Y => Delay64No3_out);

   Delay64No5_instance: Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=44 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1206_out,
                 Y => Delay64No5_out);

   Delay15No26_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg900_out,
                 Y => Delay15No26_out);

   Delay78No24_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1090_out,
                 Y => Delay78No24_out);

   Delay78No25_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg942_out,
                 Y => Delay78No25_out);

   Delay78No27_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1136_out,
                 Y => Delay78No27_out);

   Delay78No29_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1058_out,
                 Y => Delay78No29_out);

   Delay80No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1147_out,
                 Y => Delay80No_out);

   Delay80No1_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1069_out,
                 Y => Delay80No1_out);

   Delay80No2_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1027_out,
                 Y => Delay80No2_out);

   Delay80No3_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1043_out,
                 Y => Delay80No3_out);

   Delay80No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1126_out,
                 Y => Delay80No4_out);

   Delay80No5_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1114_out,
                 Y => Delay80No5_out);

   Delay87No12_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg990_out,
                 Y => Delay87No12_out);

   Delay87No13_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1001_out,
                 Y => Delay87No13_out);

   Delay87No14_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1010_out,
                 Y => Delay87No14_out);

   Delay87No15_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1103_out,
                 Y => Delay87No15_out);

   Delay87No16_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg976_out,
                 Y => Delay87No16_out);

   Delay87No17_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1254_out,
                 Y => Delay87No17_out);

   MUX_Add141_5_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add141_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Add141_5_impl_0_LUT_out);

   MUX_Add141_5_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add141_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Add141_5_impl_1_LUT_out);

   MUX_Product62_5_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product62_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Product62_5_impl_0_LUT_out);

   MUX_Product62_5_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product62_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Product62_5_impl_1_LUT_out);

   MUX_Add10_5_impl_0_LUT_instance: GenericLut_LUTData_MUX_Add10_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Add10_5_impl_0_LUT_out);

   MUX_Add10_5_impl_1_LUT_instance: GenericLut_LUTData_MUX_Add10_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Add10_5_impl_1_LUT_out);

   MUX_Divide_0_impl_0_LUT_instance: GenericLut_LUTData_MUX_Divide_0_impl_0_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Divide_0_impl_0_LUT_out);

   MUX_Divide_0_impl_1_LUT_instance: GenericLut_LUTData_MUX_Divide_0_impl_1_LUT_wIn_4_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Divide_0_impl_1_LUT_out);

   MUX_Product213_5_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product213_5_impl_0_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Product213_5_impl_0_LUT_out);

   MUX_Product213_5_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product213_5_impl_1_LUT_wIn_4_wOut_4_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount131_out,
                 Output => MUX_Product213_5_impl_1_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UV_del_1_0_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg2_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg3_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg4_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg5_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg6_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg7_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg8_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg9_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UV_del_1_1_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg11_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg12_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg13_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg14_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg15_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg16_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg17_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg18_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg19_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg20_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UV_del_1_2_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg22_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg23_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg24_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg25_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg26_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg27_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg28_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg29_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg30_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg31_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UV_del_1_3_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg33_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg34_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg35_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg36_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg37_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg38_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg39_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg40_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UV_del_1_4_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg47_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UV_del_1_5_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg55_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg63_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UW_del_1_0_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg69_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=48 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg71_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg73_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UW_del_1_1_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg76_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg80_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=48 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg81_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg82_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UW_del_1_2_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg86_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg87_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg88_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg89_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg90_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=48 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg92_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg93_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg94_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UW_del_1_3_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg97_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg98_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg99_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg100_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=48 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg101_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg102_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg103_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg104_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UW_del_1_4_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg106_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg108_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg110_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=48 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg112_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg113_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_UW_del_1_5_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg117_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg118_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=48 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg121_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg123_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VU_del_1_0_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg126_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg129_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg132_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VU_del_1_1_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg134_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg139_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg140_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VU_del_1_2_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg143_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg144_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg145_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg146_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VU_del_1_3_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg152_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg153_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg156_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VU_del_1_4_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg158_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg160_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg161_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg162_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg163_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg164_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VU_del_1_5_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg166_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg167_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg168_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg169_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg170_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg171_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg172_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VW_del_1_0_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg174_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg176_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg178_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg179_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg180_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg181_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg182_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg183_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VW_del_1_1_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg185_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg186_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg187_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg190_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg191_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg192_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg193_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg194_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VW_del_1_2_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg196_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg197_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg198_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg200_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg201_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg202_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg203_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg204_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg205_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VW_del_1_3_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg207_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg208_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg209_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg210_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg211_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg212_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg213_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg214_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg215_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg216_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VW_del_1_4_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg218_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg219_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg220_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg221_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg222_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg223_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg224_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg225_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg226_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg227_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_VW_del_1_5_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg229_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg230_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg231_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg232_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg233_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg234_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg235_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg236_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg237_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg238_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WU_del_1_0_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg240_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg241_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg242_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg243_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=42 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg244_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg245_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg246_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg247_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg248_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WU_del_1_1_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg250_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg251_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg252_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg253_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=42 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg254_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg255_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg256_out,
                 Y => SharedReg257_out);

   SharedReg258_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg257_out,
                 Y => SharedReg258_out);

   SharedReg259_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg258_out,
                 Y => SharedReg259_out);

   SharedReg260_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WU_del_1_2_out,
                 Y => SharedReg260_out);

   SharedReg261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg260_out,
                 Y => SharedReg261_out);

   SharedReg262_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg261_out,
                 Y => SharedReg262_out);

   SharedReg263_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg262_out,
                 Y => SharedReg263_out);

   SharedReg264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg263_out,
                 Y => SharedReg264_out);

   SharedReg265_instance: Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=42 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg264_out,
                 Y => SharedReg265_out);

   SharedReg266_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg265_out,
                 Y => SharedReg266_out);

   SharedReg267_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg266_out,
                 Y => SharedReg267_out);

   SharedReg268_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg267_out,
                 Y => SharedReg268_out);

   SharedReg269_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg268_out,
                 Y => SharedReg269_out);

   SharedReg270_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WU_del_1_3_out,
                 Y => SharedReg270_out);

   SharedReg271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg270_out,
                 Y => SharedReg271_out);

   SharedReg272_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg271_out,
                 Y => SharedReg272_out);

   SharedReg273_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg272_out,
                 Y => SharedReg273_out);

   SharedReg274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg273_out,
                 Y => SharedReg274_out);

   SharedReg275_instance: Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=42 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg274_out,
                 Y => SharedReg275_out);

   SharedReg276_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg275_out,
                 Y => SharedReg276_out);

   SharedReg277_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg276_out,
                 Y => SharedReg277_out);

   SharedReg278_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg277_out,
                 Y => SharedReg278_out);

   SharedReg279_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg278_out,
                 Y => SharedReg279_out);

   SharedReg280_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WU_del_1_4_out,
                 Y => SharedReg280_out);

   SharedReg281_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg280_out,
                 Y => SharedReg281_out);

   SharedReg282_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg281_out,
                 Y => SharedReg282_out);

   SharedReg283_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg282_out,
                 Y => SharedReg283_out);

   SharedReg284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg283_out,
                 Y => SharedReg284_out);

   SharedReg285_instance: Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=42 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg284_out,
                 Y => SharedReg285_out);

   SharedReg286_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg285_out,
                 Y => SharedReg286_out);

   SharedReg287_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg286_out,
                 Y => SharedReg287_out);

   SharedReg288_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg287_out,
                 Y => SharedReg288_out);

   SharedReg289_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg288_out,
                 Y => SharedReg289_out);

   SharedReg290_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WU_del_1_5_out,
                 Y => SharedReg290_out);

   SharedReg291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg290_out,
                 Y => SharedReg291_out);

   SharedReg292_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg291_out,
                 Y => SharedReg292_out);

   SharedReg293_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg292_out,
                 Y => SharedReg293_out);

   SharedReg294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg293_out,
                 Y => SharedReg294_out);

   SharedReg295_instance: Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=42 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg294_out,
                 Y => SharedReg295_out);

   SharedReg296_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg295_out,
                 Y => SharedReg296_out);

   SharedReg297_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg296_out,
                 Y => SharedReg297_out);

   SharedReg298_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg297_out,
                 Y => SharedReg298_out);

   SharedReg299_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg298_out,
                 Y => SharedReg299_out);

   SharedReg300_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WV_del_1_0_out,
                 Y => SharedReg300_out);

   SharedReg301_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg300_out,
                 Y => SharedReg301_out);

   SharedReg302_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg301_out,
                 Y => SharedReg302_out);

   SharedReg303_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg302_out,
                 Y => SharedReg303_out);

   SharedReg304_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg303_out,
                 Y => SharedReg304_out);

   SharedReg305_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg304_out,
                 Y => SharedReg305_out);

   SharedReg306_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg305_out,
                 Y => SharedReg306_out);

   SharedReg307_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg306_out,
                 Y => SharedReg307_out);

   SharedReg308_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg307_out,
                 Y => SharedReg308_out);

   SharedReg309_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WV_del_1_1_out,
                 Y => SharedReg309_out);

   SharedReg310_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg309_out,
                 Y => SharedReg310_out);

   SharedReg311_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg310_out,
                 Y => SharedReg311_out);

   SharedReg312_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg311_out,
                 Y => SharedReg312_out);

   SharedReg313_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg312_out,
                 Y => SharedReg313_out);

   SharedReg314_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg313_out,
                 Y => SharedReg314_out);

   SharedReg315_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg314_out,
                 Y => SharedReg315_out);

   SharedReg316_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg315_out,
                 Y => SharedReg316_out);

   SharedReg317_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg316_out,
                 Y => SharedReg317_out);

   SharedReg318_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WV_del_1_2_out,
                 Y => SharedReg318_out);

   SharedReg319_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg318_out,
                 Y => SharedReg319_out);

   SharedReg320_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg319_out,
                 Y => SharedReg320_out);

   SharedReg321_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg320_out,
                 Y => SharedReg321_out);

   SharedReg322_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg321_out,
                 Y => SharedReg322_out);

   SharedReg323_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg322_out,
                 Y => SharedReg323_out);

   SharedReg324_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg323_out,
                 Y => SharedReg324_out);

   SharedReg325_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg324_out,
                 Y => SharedReg325_out);

   SharedReg326_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg325_out,
                 Y => SharedReg326_out);

   SharedReg327_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WV_del_1_3_out,
                 Y => SharedReg327_out);

   SharedReg328_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg327_out,
                 Y => SharedReg328_out);

   SharedReg329_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg328_out,
                 Y => SharedReg329_out);

   SharedReg330_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg329_out,
                 Y => SharedReg330_out);

   SharedReg331_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg330_out,
                 Y => SharedReg331_out);

   SharedReg332_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg331_out,
                 Y => SharedReg332_out);

   SharedReg333_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg332_out,
                 Y => SharedReg333_out);

   SharedReg334_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg333_out,
                 Y => SharedReg334_out);

   SharedReg335_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg334_out,
                 Y => SharedReg335_out);

   SharedReg336_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WV_del_1_4_out,
                 Y => SharedReg336_out);

   SharedReg337_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg336_out,
                 Y => SharedReg337_out);

   SharedReg338_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg337_out,
                 Y => SharedReg338_out);

   SharedReg339_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg338_out,
                 Y => SharedReg339_out);

   SharedReg340_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg339_out,
                 Y => SharedReg340_out);

   SharedReg341_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg340_out,
                 Y => SharedReg341_out);

   SharedReg342_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg341_out,
                 Y => SharedReg342_out);

   SharedReg343_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg342_out,
                 Y => SharedReg343_out);

   SharedReg344_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg343_out,
                 Y => SharedReg344_out);

   SharedReg345_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Ldiff_WV_del_1_5_out,
                 Y => SharedReg345_out);

   SharedReg346_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg345_out,
                 Y => SharedReg346_out);

   SharedReg347_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg346_out,
                 Y => SharedReg347_out);

   SharedReg348_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg347_out,
                 Y => SharedReg348_out);

   SharedReg349_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg348_out,
                 Y => SharedReg349_out);

   SharedReg350_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg349_out,
                 Y => SharedReg350_out);

   SharedReg351_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg350_out,
                 Y => SharedReg351_out);

   SharedReg352_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg351_out,
                 Y => SharedReg352_out);

   SharedReg353_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg352_out,
                 Y => SharedReg353_out);

   SharedReg354_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_0_impl_out,
                 Y => SharedReg354_out);

   SharedReg355_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg354_out,
                 Y => SharedReg355_out);

   SharedReg356_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg355_out,
                 Y => SharedReg356_out);

   SharedReg357_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg356_out,
                 Y => SharedReg357_out);

   SharedReg358_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg357_out,
                 Y => SharedReg358_out);

   SharedReg359_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg358_out,
                 Y => SharedReg359_out);

   SharedReg360_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg359_out,
                 Y => SharedReg360_out);

   SharedReg361_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg360_out,
                 Y => SharedReg361_out);

   SharedReg362_instance: Delay_34_DelayLength_78_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=78 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg361_out,
                 Y => SharedReg362_out);

   SharedReg363_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_1_impl_out,
                 Y => SharedReg363_out);

   SharedReg364_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg363_out,
                 Y => SharedReg364_out);

   SharedReg365_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg364_out,
                 Y => SharedReg365_out);

   SharedReg366_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg365_out,
                 Y => SharedReg366_out);

   SharedReg367_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg366_out,
                 Y => SharedReg367_out);

   SharedReg368_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg367_out,
                 Y => SharedReg368_out);

   SharedReg369_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg368_out,
                 Y => SharedReg369_out);

   SharedReg370_instance: Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=67 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg369_out,
                 Y => SharedReg370_out);

   SharedReg371_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_2_impl_out,
                 Y => SharedReg371_out);

   SharedReg372_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg371_out,
                 Y => SharedReg372_out);

   SharedReg373_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg372_out,
                 Y => SharedReg373_out);

   SharedReg374_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg373_out,
                 Y => SharedReg374_out);

   SharedReg375_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg374_out,
                 Y => SharedReg375_out);

   SharedReg376_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg375_out,
                 Y => SharedReg376_out);

   SharedReg377_instance: Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=38 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg376_out,
                 Y => SharedReg377_out);

   SharedReg378_instance: Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=39 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg377_out,
                 Y => SharedReg378_out);

   SharedReg379_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_3_impl_out,
                 Y => SharedReg379_out);

   SharedReg380_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg379_out,
                 Y => SharedReg380_out);

   SharedReg381_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg380_out,
                 Y => SharedReg381_out);

   SharedReg382_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg381_out,
                 Y => SharedReg382_out);

   SharedReg383_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg382_out,
                 Y => SharedReg383_out);

   SharedReg384_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg383_out,
                 Y => SharedReg384_out);

   SharedReg385_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg384_out,
                 Y => SharedReg385_out);

   SharedReg386_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_4_impl_out,
                 Y => SharedReg386_out);

   SharedReg387_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg386_out,
                 Y => SharedReg387_out);

   SharedReg388_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg387_out,
                 Y => SharedReg388_out);

   SharedReg389_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg388_out,
                 Y => SharedReg389_out);

   SharedReg390_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg389_out,
                 Y => SharedReg390_out);

   SharedReg391_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg390_out,
                 Y => SharedReg391_out);

   SharedReg392_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg391_out,
                 Y => SharedReg392_out);

   SharedReg393_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg392_out,
                 Y => SharedReg393_out);

   SharedReg394_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product108_5_impl_out,
                 Y => SharedReg394_out);

   SharedReg395_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg394_out,
                 Y => SharedReg395_out);

   SharedReg396_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg395_out,
                 Y => SharedReg396_out);

   SharedReg397_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg396_out,
                 Y => SharedReg397_out);

   SharedReg398_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg397_out,
                 Y => SharedReg398_out);

   SharedReg399_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg398_out,
                 Y => SharedReg399_out);

   SharedReg400_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_0_impl_out,
                 Y => SharedReg400_out);

   SharedReg401_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg400_out,
                 Y => SharedReg401_out);

   SharedReg402_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg401_out,
                 Y => SharedReg402_out);

   SharedReg403_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg402_out,
                 Y => SharedReg403_out);

   SharedReg404_instance: Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=55 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg403_out,
                 Y => SharedReg404_out);

   SharedReg405_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg404_out,
                 Y => SharedReg405_out);

   SharedReg406_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg405_out,
                 Y => SharedReg406_out);

   SharedReg407_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg406_out,
                 Y => SharedReg407_out);

   SharedReg408_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_1_impl_out,
                 Y => SharedReg408_out);

   SharedReg409_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg408_out,
                 Y => SharedReg409_out);

   SharedReg410_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg409_out,
                 Y => SharedReg410_out);

   SharedReg411_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg410_out,
                 Y => SharedReg411_out);

   SharedReg412_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg411_out,
                 Y => SharedReg412_out);

   SharedReg413_instance: Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=53 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg412_out,
                 Y => SharedReg413_out);

   SharedReg414_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg413_out,
                 Y => SharedReg414_out);

   SharedReg415_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg414_out,
                 Y => SharedReg415_out);

   SharedReg416_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg415_out,
                 Y => SharedReg416_out);

   SharedReg417_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg416_out,
                 Y => SharedReg417_out);

   SharedReg418_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_2_impl_out,
                 Y => SharedReg418_out);

   SharedReg419_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg418_out,
                 Y => SharedReg419_out);

   SharedReg420_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg419_out,
                 Y => SharedReg420_out);

   SharedReg421_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg420_out,
                 Y => SharedReg421_out);

   SharedReg422_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg421_out,
                 Y => SharedReg422_out);

   SharedReg423_instance: Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=53 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg422_out,
                 Y => SharedReg423_out);

   SharedReg424_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg423_out,
                 Y => SharedReg424_out);

   SharedReg425_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_3_impl_out,
                 Y => SharedReg425_out);

   SharedReg426_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg425_out,
                 Y => SharedReg426_out);

   SharedReg427_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg426_out,
                 Y => SharedReg427_out);

   SharedReg428_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg427_out,
                 Y => SharedReg428_out);

   SharedReg429_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg428_out,
                 Y => SharedReg429_out);

   SharedReg430_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg429_out,
                 Y => SharedReg430_out);

   SharedReg431_instance: Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=55 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg430_out,
                 Y => SharedReg431_out);

   SharedReg432_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg431_out,
                 Y => SharedReg432_out);

   SharedReg433_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_4_impl_out,
                 Y => SharedReg433_out);

   SharedReg434_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg433_out,
                 Y => SharedReg434_out);

   SharedReg435_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg434_out,
                 Y => SharedReg435_out);

   SharedReg436_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg435_out,
                 Y => SharedReg436_out);

   SharedReg437_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg436_out,
                 Y => SharedReg437_out);

   SharedReg438_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg437_out,
                 Y => SharedReg438_out);

   SharedReg439_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg438_out,
                 Y => SharedReg439_out);

   SharedReg440_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg439_out,
                 Y => SharedReg440_out);

   SharedReg441_instance: Delay_34_DelayLength_55_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=55 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg440_out,
                 Y => SharedReg441_out);

   SharedReg442_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product110_5_impl_out,
                 Y => SharedReg442_out);

   SharedReg443_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg442_out,
                 Y => SharedReg443_out);

   SharedReg444_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg443_out,
                 Y => SharedReg444_out);

   SharedReg445_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg444_out,
                 Y => SharedReg445_out);

   SharedReg446_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg445_out,
                 Y => SharedReg446_out);

   SharedReg447_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg446_out,
                 Y => SharedReg447_out);

   SharedReg448_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg447_out,
                 Y => SharedReg448_out);

   SharedReg449_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg448_out,
                 Y => SharedReg449_out);

   SharedReg450_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product109_0_impl_out,
                 Y => SharedReg450_out);

   SharedReg451_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg450_out,
                 Y => SharedReg451_out);

   SharedReg452_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg451_out,
                 Y => SharedReg452_out);

   SharedReg453_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg452_out,
                 Y => SharedReg453_out);

   SharedReg454_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg453_out,
                 Y => SharedReg454_out);

   SharedReg455_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg454_out,
                 Y => SharedReg455_out);

   SharedReg456_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product109_1_impl_out,
                 Y => SharedReg456_out);

   SharedReg457_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg456_out,
                 Y => SharedReg457_out);

   SharedReg458_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg457_out,
                 Y => SharedReg458_out);

   SharedReg459_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg458_out,
                 Y => SharedReg459_out);

   SharedReg460_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg459_out,
                 Y => SharedReg460_out);

   SharedReg461_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg460_out,
                 Y => SharedReg461_out);

   SharedReg462_instance: Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=42 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg461_out,
                 Y => SharedReg462_out);

   SharedReg463_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product109_2_impl_out,
                 Y => SharedReg463_out);

   SharedReg464_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg463_out,
                 Y => SharedReg464_out);

   SharedReg465_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg464_out,
                 Y => SharedReg465_out);

   SharedReg466_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg465_out,
                 Y => SharedReg466_out);

   SharedReg467_instance: Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=42 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg466_out,
                 Y => SharedReg467_out);

   SharedReg468_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg467_out,
                 Y => SharedReg468_out);

   SharedReg469_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg468_out,
                 Y => SharedReg469_out);

   SharedReg470_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg469_out,
                 Y => SharedReg470_out);

   SharedReg471_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product109_3_impl_out,
                 Y => SharedReg471_out);

   SharedReg472_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg471_out,
                 Y => SharedReg472_out);

   SharedReg473_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg472_out,
                 Y => SharedReg473_out);

   SharedReg474_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg473_out,
                 Y => SharedReg474_out);

   SharedReg475_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg474_out,
                 Y => SharedReg475_out);

   SharedReg476_instance: Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=47 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg475_out,
                 Y => SharedReg476_out);

   SharedReg477_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg476_out,
                 Y => SharedReg477_out);

   SharedReg478_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg477_out,
                 Y => SharedReg478_out);

   SharedReg479_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product109_4_impl_out,
                 Y => SharedReg479_out);

   SharedReg480_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg479_out,
                 Y => SharedReg480_out);

   SharedReg481_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg480_out,
                 Y => SharedReg481_out);

   SharedReg482_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg481_out,
                 Y => SharedReg482_out);

   SharedReg483_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg482_out,
                 Y => SharedReg483_out);

   SharedReg484_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg483_out,
                 Y => SharedReg484_out);

   SharedReg485_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg484_out,
                 Y => SharedReg485_out);

   SharedReg486_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg485_out,
                 Y => SharedReg486_out);

   SharedReg487_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product109_5_impl_out,
                 Y => SharedReg487_out);

   SharedReg488_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg487_out,
                 Y => SharedReg488_out);

   SharedReg489_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg488_out,
                 Y => SharedReg489_out);

   SharedReg490_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg489_out,
                 Y => SharedReg490_out);

   SharedReg491_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg490_out,
                 Y => SharedReg491_out);

   SharedReg492_instance: Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=43 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg491_out,
                 Y => SharedReg492_out);

   SharedReg493_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_0_impl_out,
                 Y => SharedReg493_out);

   SharedReg494_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg493_out,
                 Y => SharedReg494_out);

   SharedReg495_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg494_out,
                 Y => SharedReg495_out);

   SharedReg496_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg495_out,
                 Y => SharedReg496_out);

   SharedReg497_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg496_out,
                 Y => SharedReg497_out);

   SharedReg498_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg497_out,
                 Y => SharedReg498_out);

   SharedReg499_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_1_impl_out,
                 Y => SharedReg499_out);

   SharedReg500_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg499_out,
                 Y => SharedReg500_out);

   SharedReg501_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg500_out,
                 Y => SharedReg501_out);

   SharedReg502_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg501_out,
                 Y => SharedReg502_out);

   SharedReg503_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg502_out,
                 Y => SharedReg503_out);

   SharedReg504_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_2_impl_out,
                 Y => SharedReg504_out);

   SharedReg505_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg504_out,
                 Y => SharedReg505_out);

   SharedReg506_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg505_out,
                 Y => SharedReg506_out);

   SharedReg507_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg506_out,
                 Y => SharedReg507_out);

   SharedReg508_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg507_out,
                 Y => SharedReg508_out);

   SharedReg509_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg508_out,
                 Y => SharedReg509_out);

   SharedReg510_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg509_out,
                 Y => SharedReg510_out);

   SharedReg511_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_3_impl_out,
                 Y => SharedReg511_out);

   SharedReg512_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg511_out,
                 Y => SharedReg512_out);

   SharedReg513_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg512_out,
                 Y => SharedReg513_out);

   SharedReg514_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg513_out,
                 Y => SharedReg514_out);

   SharedReg515_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg514_out,
                 Y => SharedReg515_out);

   SharedReg516_instance: Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=47 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg515_out,
                 Y => SharedReg516_out);

   SharedReg517_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_4_impl_out,
                 Y => SharedReg517_out);

   SharedReg518_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg517_out,
                 Y => SharedReg518_out);

   SharedReg519_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg518_out,
                 Y => SharedReg519_out);

   SharedReg520_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg519_out,
                 Y => SharedReg520_out);

   SharedReg521_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg520_out,
                 Y => SharedReg521_out);

   SharedReg522_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg521_out,
                 Y => SharedReg522_out);

   SharedReg523_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg522_out,
                 Y => SharedReg523_out);

   SharedReg524_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product111_5_impl_out,
                 Y => SharedReg524_out);

   SharedReg525_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg524_out,
                 Y => SharedReg525_out);

   SharedReg526_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg525_out,
                 Y => SharedReg526_out);

   SharedReg527_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg526_out,
                 Y => SharedReg527_out);

   SharedReg528_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg527_out,
                 Y => SharedReg528_out);

   SharedReg529_instance: Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=63 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg528_out,
                 Y => SharedReg529_out);

   SharedReg530_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg529_out,
                 Y => SharedReg530_out);

   SharedReg531_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_0_impl_out,
                 Y => SharedReg531_out);

   SharedReg532_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg531_out,
                 Y => SharedReg532_out);

   SharedReg533_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg532_out,
                 Y => SharedReg533_out);

   SharedReg534_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg533_out,
                 Y => SharedReg534_out);

   SharedReg535_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg534_out,
                 Y => SharedReg535_out);

   SharedReg536_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg535_out,
                 Y => SharedReg536_out);

   SharedReg537_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg536_out,
                 Y => SharedReg537_out);

   SharedReg538_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg537_out,
                 Y => SharedReg538_out);

   SharedReg539_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg538_out,
                 Y => SharedReg539_out);

   SharedReg540_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_1_impl_out,
                 Y => SharedReg540_out);

   SharedReg541_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg540_out,
                 Y => SharedReg541_out);

   SharedReg542_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg541_out,
                 Y => SharedReg542_out);

   SharedReg543_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg542_out,
                 Y => SharedReg543_out);

   SharedReg544_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg543_out,
                 Y => SharedReg544_out);

   SharedReg545_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg544_out,
                 Y => SharedReg545_out);

   SharedReg546_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg545_out,
                 Y => SharedReg546_out);

   SharedReg547_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg546_out,
                 Y => SharedReg547_out);

   SharedReg548_instance: Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=58 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg547_out,
                 Y => SharedReg548_out);

   SharedReg549_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg548_out,
                 Y => SharedReg549_out);

   SharedReg550_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_2_impl_out,
                 Y => SharedReg550_out);

   SharedReg551_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg550_out,
                 Y => SharedReg551_out);

   SharedReg552_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg551_out,
                 Y => SharedReg552_out);

   SharedReg553_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg552_out,
                 Y => SharedReg553_out);

   SharedReg554_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg553_out,
                 Y => SharedReg554_out);

   SharedReg555_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg554_out,
                 Y => SharedReg555_out);

   SharedReg556_instance: Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=62 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg555_out,
                 Y => SharedReg556_out);

   SharedReg557_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_3_impl_out,
                 Y => SharedReg557_out);

   SharedReg558_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg557_out,
                 Y => SharedReg558_out);

   SharedReg559_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg558_out,
                 Y => SharedReg559_out);

   SharedReg560_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg559_out,
                 Y => SharedReg560_out);

   SharedReg561_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg560_out,
                 Y => SharedReg561_out);

   SharedReg562_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg561_out,
                 Y => SharedReg562_out);

   SharedReg563_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg562_out,
                 Y => SharedReg563_out);

   SharedReg564_instance: Delay_34_DelayLength_51_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=51 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg563_out,
                 Y => SharedReg564_out);

   SharedReg565_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg564_out,
                 Y => SharedReg565_out);

   SharedReg566_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_4_impl_out,
                 Y => SharedReg566_out);

   SharedReg567_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg566_out,
                 Y => SharedReg567_out);

   SharedReg568_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg567_out,
                 Y => SharedReg568_out);

   SharedReg569_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg568_out,
                 Y => SharedReg569_out);

   SharedReg570_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg569_out,
                 Y => SharedReg570_out);

   SharedReg571_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg570_out,
                 Y => SharedReg571_out);

   SharedReg572_instance: Delay_34_DelayLength_63_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=63 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg571_out,
                 Y => SharedReg572_out);

   SharedReg573_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product210_5_impl_out,
                 Y => SharedReg573_out);

   SharedReg574_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg573_out,
                 Y => SharedReg574_out);

   SharedReg575_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg574_out,
                 Y => SharedReg575_out);

   SharedReg576_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg575_out,
                 Y => SharedReg576_out);

   SharedReg577_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg576_out,
                 Y => SharedReg577_out);

   SharedReg578_instance: Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=48 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg577_out,
                 Y => SharedReg578_out);

   SharedReg579_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg578_out,
                 Y => SharedReg579_out);

   SharedReg580_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg579_out,
                 Y => SharedReg580_out);

   SharedReg581_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_0_impl_out,
                 Y => SharedReg581_out);

   SharedReg582_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg581_out,
                 Y => SharedReg582_out);

   SharedReg583_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg582_out,
                 Y => SharedReg583_out);

   SharedReg584_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg583_out,
                 Y => SharedReg584_out);

   SharedReg585_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg584_out,
                 Y => SharedReg585_out);

   SharedReg586_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg585_out,
                 Y => SharedReg586_out);

   SharedReg587_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg586_out,
                 Y => SharedReg587_out);

   SharedReg588_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg587_out,
                 Y => SharedReg588_out);

   SharedReg589_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_1_impl_out,
                 Y => SharedReg589_out);

   SharedReg590_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg589_out,
                 Y => SharedReg590_out);

   SharedReg591_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg590_out,
                 Y => SharedReg591_out);

   SharedReg592_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg591_out,
                 Y => SharedReg592_out);

   SharedReg593_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg592_out,
                 Y => SharedReg593_out);

   SharedReg594_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg593_out,
                 Y => SharedReg594_out);

   SharedReg595_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg594_out,
                 Y => SharedReg595_out);

   SharedReg596_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg595_out,
                 Y => SharedReg596_out);

   SharedReg597_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_2_impl_out,
                 Y => SharedReg597_out);

   SharedReg598_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg597_out,
                 Y => SharedReg598_out);

   SharedReg599_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg598_out,
                 Y => SharedReg599_out);

   SharedReg600_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg599_out,
                 Y => SharedReg600_out);

   SharedReg601_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg600_out,
                 Y => SharedReg601_out);

   SharedReg602_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg601_out,
                 Y => SharedReg602_out);

   SharedReg603_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg602_out,
                 Y => SharedReg603_out);

   SharedReg604_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg603_out,
                 Y => SharedReg604_out);

   SharedReg605_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_3_impl_out,
                 Y => SharedReg605_out);

   SharedReg606_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg605_out,
                 Y => SharedReg606_out);

   SharedReg607_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg606_out,
                 Y => SharedReg607_out);

   SharedReg608_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg607_out,
                 Y => SharedReg608_out);

   SharedReg609_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg608_out,
                 Y => SharedReg609_out);

   SharedReg610_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_4_impl_out,
                 Y => SharedReg610_out);

   SharedReg611_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg610_out,
                 Y => SharedReg611_out);

   SharedReg612_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg611_out,
                 Y => SharedReg612_out);

   SharedReg613_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg612_out,
                 Y => SharedReg613_out);

   SharedReg614_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg613_out,
                 Y => SharedReg614_out);

   SharedReg615_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg614_out,
                 Y => SharedReg615_out);

   SharedReg616_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg615_out,
                 Y => SharedReg616_out);

   SharedReg617_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg616_out,
                 Y => SharedReg617_out);

   SharedReg618_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product310_5_impl_out,
                 Y => SharedReg618_out);

   SharedReg619_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg618_out,
                 Y => SharedReg619_out);

   SharedReg620_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg619_out,
                 Y => SharedReg620_out);

   SharedReg621_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg620_out,
                 Y => SharedReg621_out);

   SharedReg622_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg621_out,
                 Y => SharedReg622_out);

   SharedReg623_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg622_out,
                 Y => SharedReg623_out);

   SharedReg624_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg623_out,
                 Y => SharedReg624_out);

   SharedReg625_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg624_out,
                 Y => SharedReg625_out);

   SharedReg626_instance: Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=42 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg625_out,
                 Y => SharedReg626_out);

   SharedReg627_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product410_0_impl_out,
                 Y => SharedReg627_out);

   SharedReg628_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg627_out,
                 Y => SharedReg628_out);

   SharedReg629_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg628_out,
                 Y => SharedReg629_out);

   SharedReg630_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg629_out,
                 Y => SharedReg630_out);

   SharedReg631_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg630_out,
                 Y => SharedReg631_out);

   SharedReg632_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg631_out,
                 Y => SharedReg632_out);

   SharedReg633_instance: Delay_34_DelayLength_46_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=46 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg632_out,
                 Y => SharedReg633_out);

   SharedReg634_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product410_1_impl_out,
                 Y => SharedReg634_out);

   SharedReg635_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg634_out,
                 Y => SharedReg635_out);

   SharedReg636_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg635_out,
                 Y => SharedReg636_out);

   SharedReg637_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg636_out,
                 Y => SharedReg637_out);

   SharedReg638_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg637_out,
                 Y => SharedReg638_out);

   SharedReg639_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg638_out,
                 Y => SharedReg639_out);

   SharedReg640_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg639_out,
                 Y => SharedReg640_out);

   SharedReg641_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg640_out,
                 Y => SharedReg641_out);

   SharedReg642_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product410_2_impl_out,
                 Y => SharedReg642_out);

   SharedReg643_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg642_out,
                 Y => SharedReg643_out);

   SharedReg644_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg643_out,
                 Y => SharedReg644_out);

   SharedReg645_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg644_out,
                 Y => SharedReg645_out);

   SharedReg646_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg645_out,
                 Y => SharedReg646_out);

   SharedReg647_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg646_out,
                 Y => SharedReg647_out);

   SharedReg648_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg647_out,
                 Y => SharedReg648_out);

   SharedReg649_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg648_out,
                 Y => SharedReg649_out);

   SharedReg650_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg649_out,
                 Y => SharedReg650_out);

   SharedReg651_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg650_out,
                 Y => SharedReg651_out);

   SharedReg652_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product410_3_impl_out,
                 Y => SharedReg652_out);

   SharedReg653_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg652_out,
                 Y => SharedReg653_out);

   SharedReg654_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg653_out,
                 Y => SharedReg654_out);

   SharedReg655_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg654_out,
                 Y => SharedReg655_out);

   SharedReg656_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg655_out,
                 Y => SharedReg656_out);

   SharedReg657_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg656_out,
                 Y => SharedReg657_out);

   SharedReg658_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg657_out,
                 Y => SharedReg658_out);

   SharedReg659_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg658_out,
                 Y => SharedReg659_out);

   SharedReg660_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg659_out,
                 Y => SharedReg660_out);

   SharedReg661_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product410_4_impl_out,
                 Y => SharedReg661_out);

   SharedReg662_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg661_out,
                 Y => SharedReg662_out);

   SharedReg663_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg662_out,
                 Y => SharedReg663_out);

   SharedReg664_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg663_out,
                 Y => SharedReg664_out);

   SharedReg665_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg664_out,
                 Y => SharedReg665_out);

   SharedReg666_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg665_out,
                 Y => SharedReg666_out);

   SharedReg667_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg666_out,
                 Y => SharedReg667_out);

   SharedReg668_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg667_out,
                 Y => SharedReg668_out);

   SharedReg669_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product410_5_impl_out,
                 Y => SharedReg669_out);

   SharedReg670_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg669_out,
                 Y => SharedReg670_out);

   SharedReg671_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg670_out,
                 Y => SharedReg671_out);

   SharedReg672_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg671_out,
                 Y => SharedReg672_out);

   SharedReg673_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg672_out,
                 Y => SharedReg673_out);

   SharedReg674_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg673_out,
                 Y => SharedReg674_out);

   SharedReg675_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg674_out,
                 Y => SharedReg675_out);

   SharedReg676_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product510_0_impl_out,
                 Y => SharedReg676_out);

   SharedReg677_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg676_out,
                 Y => SharedReg677_out);

   SharedReg678_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg677_out,
                 Y => SharedReg678_out);

   SharedReg679_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg678_out,
                 Y => SharedReg679_out);

   SharedReg680_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg679_out,
                 Y => SharedReg680_out);

   SharedReg681_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg680_out,
                 Y => SharedReg681_out);

   SharedReg682_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg681_out,
                 Y => SharedReg682_out);

   SharedReg683_instance: Delay_34_DelayLength_53_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=53 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg682_out,
                 Y => SharedReg683_out);

   SharedReg684_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product510_1_impl_out,
                 Y => SharedReg684_out);

   SharedReg685_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg684_out,
                 Y => SharedReg685_out);

   SharedReg686_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg685_out,
                 Y => SharedReg686_out);

   SharedReg687_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg686_out,
                 Y => SharedReg687_out);

   SharedReg688_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg687_out,
                 Y => SharedReg688_out);

   SharedReg689_instance: Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=62 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg688_out,
                 Y => SharedReg689_out);

   SharedReg690_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product510_2_impl_out,
                 Y => SharedReg690_out);

   SharedReg691_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg690_out,
                 Y => SharedReg691_out);

   SharedReg692_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg691_out,
                 Y => SharedReg692_out);

   SharedReg693_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg692_out,
                 Y => SharedReg693_out);

   SharedReg694_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg693_out,
                 Y => SharedReg694_out);

   SharedReg695_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg694_out,
                 Y => SharedReg695_out);

   SharedReg696_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg695_out,
                 Y => SharedReg696_out);

   SharedReg697_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg696_out,
                 Y => SharedReg697_out);

   SharedReg698_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg697_out,
                 Y => SharedReg698_out);

   SharedReg699_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg698_out,
                 Y => SharedReg699_out);

   SharedReg700_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product510_3_impl_out,
                 Y => SharedReg700_out);

   SharedReg701_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg700_out,
                 Y => SharedReg701_out);

   SharedReg702_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg701_out,
                 Y => SharedReg702_out);

   SharedReg703_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg702_out,
                 Y => SharedReg703_out);

   SharedReg704_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg703_out,
                 Y => SharedReg704_out);

   SharedReg705_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg704_out,
                 Y => SharedReg705_out);

   SharedReg706_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg705_out,
                 Y => SharedReg706_out);

   SharedReg707_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg706_out,
                 Y => SharedReg707_out);

   SharedReg708_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg707_out,
                 Y => SharedReg708_out);

   SharedReg709_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product510_4_impl_out,
                 Y => SharedReg709_out);

   SharedReg710_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg709_out,
                 Y => SharedReg710_out);

   SharedReg711_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg710_out,
                 Y => SharedReg711_out);

   SharedReg712_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg711_out,
                 Y => SharedReg712_out);

   SharedReg713_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg712_out,
                 Y => SharedReg713_out);

   SharedReg714_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg713_out,
                 Y => SharedReg714_out);

   SharedReg715_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg714_out,
                 Y => SharedReg715_out);

   SharedReg716_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg715_out,
                 Y => SharedReg716_out);

   SharedReg717_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg716_out,
                 Y => SharedReg717_out);

   SharedReg718_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product510_5_impl_out,
                 Y => SharedReg718_out);

   SharedReg719_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg718_out,
                 Y => SharedReg719_out);

   SharedReg720_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg719_out,
                 Y => SharedReg720_out);

   SharedReg721_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg720_out,
                 Y => SharedReg721_out);

   SharedReg722_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg721_out,
                 Y => SharedReg722_out);

   SharedReg723_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg722_out,
                 Y => SharedReg723_out);

   SharedReg724_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg723_out,
                 Y => SharedReg724_out);

   SharedReg725_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg724_out,
                 Y => SharedReg725_out);

   SharedReg726_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_0_impl_out,
                 Y => SharedReg726_out);

   SharedReg727_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg726_out,
                 Y => SharedReg727_out);

   SharedReg728_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg727_out,
                 Y => SharedReg728_out);

   SharedReg729_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg728_out,
                 Y => SharedReg729_out);

   SharedReg730_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg729_out,
                 Y => SharedReg730_out);

   SharedReg731_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg730_out,
                 Y => SharedReg731_out);

   SharedReg732_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg731_out,
                 Y => SharedReg732_out);

   SharedReg733_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg732_out,
                 Y => SharedReg733_out);

   SharedReg734_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg733_out,
                 Y => SharedReg734_out);

   SharedReg735_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_1_impl_out,
                 Y => SharedReg735_out);

   SharedReg736_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg735_out,
                 Y => SharedReg736_out);

   SharedReg737_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg736_out,
                 Y => SharedReg737_out);

   SharedReg738_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg737_out,
                 Y => SharedReg738_out);

   SharedReg739_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg738_out,
                 Y => SharedReg739_out);

   SharedReg740_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg739_out,
                 Y => SharedReg740_out);

   SharedReg741_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg740_out,
                 Y => SharedReg741_out);

   SharedReg742_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg741_out,
                 Y => SharedReg742_out);

   SharedReg743_instance: Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=32 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg742_out,
                 Y => SharedReg743_out);

   SharedReg744_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg743_out,
                 Y => SharedReg744_out);

   SharedReg745_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg744_out,
                 Y => SharedReg745_out);

   SharedReg746_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_2_impl_out,
                 Y => SharedReg746_out);

   SharedReg747_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg746_out,
                 Y => SharedReg747_out);

   SharedReg748_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg747_out,
                 Y => SharedReg748_out);

   SharedReg749_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg748_out,
                 Y => SharedReg749_out);

   SharedReg750_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg749_out,
                 Y => SharedReg750_out);

   SharedReg751_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg750_out,
                 Y => SharedReg751_out);

   SharedReg752_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg751_out,
                 Y => SharedReg752_out);

   SharedReg753_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg752_out,
                 Y => SharedReg753_out);

   SharedReg754_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg753_out,
                 Y => SharedReg754_out);

   SharedReg755_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_3_impl_out,
                 Y => SharedReg755_out);

   SharedReg756_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg755_out,
                 Y => SharedReg756_out);

   SharedReg757_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg756_out,
                 Y => SharedReg757_out);

   SharedReg758_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg757_out,
                 Y => SharedReg758_out);

   SharedReg759_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg758_out,
                 Y => SharedReg759_out);

   SharedReg760_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg759_out,
                 Y => SharedReg760_out);

   SharedReg761_instance: Delay_34_DelayLength_48_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=48 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg760_out,
                 Y => SharedReg761_out);

   SharedReg762_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_4_impl_out,
                 Y => SharedReg762_out);

   SharedReg763_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg762_out,
                 Y => SharedReg763_out);

   SharedReg764_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg763_out,
                 Y => SharedReg764_out);

   SharedReg765_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg764_out,
                 Y => SharedReg765_out);

   SharedReg766_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg765_out,
                 Y => SharedReg766_out);

   SharedReg767_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg766_out,
                 Y => SharedReg767_out);

   SharedReg768_instance: Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=50 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg767_out,
                 Y => SharedReg768_out);

   SharedReg769_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product610_5_impl_out,
                 Y => SharedReg769_out);

   SharedReg770_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg769_out,
                 Y => SharedReg770_out);

   SharedReg771_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg770_out,
                 Y => SharedReg771_out);

   SharedReg772_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg771_out,
                 Y => SharedReg772_out);

   SharedReg773_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg772_out,
                 Y => SharedReg773_out);

   SharedReg774_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg773_out,
                 Y => SharedReg774_out);

   SharedReg775_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product710_0_impl_out,
                 Y => SharedReg775_out);

   SharedReg776_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg775_out,
                 Y => SharedReg776_out);

   SharedReg777_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg776_out,
                 Y => SharedReg777_out);

   SharedReg778_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg777_out,
                 Y => SharedReg778_out);

   SharedReg779_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg778_out,
                 Y => SharedReg779_out);

   SharedReg780_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg779_out,
                 Y => SharedReg780_out);

   SharedReg781_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg780_out,
                 Y => SharedReg781_out);

   SharedReg782_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product710_1_impl_out,
                 Y => SharedReg782_out);

   SharedReg783_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg782_out,
                 Y => SharedReg783_out);

   SharedReg784_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg783_out,
                 Y => SharedReg784_out);

   SharedReg785_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg784_out,
                 Y => SharedReg785_out);

   SharedReg786_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg785_out,
                 Y => SharedReg786_out);

   SharedReg787_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg786_out,
                 Y => SharedReg787_out);

   SharedReg788_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg787_out,
                 Y => SharedReg788_out);

   SharedReg789_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg788_out,
                 Y => SharedReg789_out);

   SharedReg790_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg789_out,
                 Y => SharedReg790_out);

   SharedReg791_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product710_2_impl_out,
                 Y => SharedReg791_out);

   SharedReg792_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg791_out,
                 Y => SharedReg792_out);

   SharedReg793_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg792_out,
                 Y => SharedReg793_out);

   SharedReg794_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg793_out,
                 Y => SharedReg794_out);

   SharedReg795_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg794_out,
                 Y => SharedReg795_out);

   SharedReg796_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg795_out,
                 Y => SharedReg796_out);

   SharedReg797_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg796_out,
                 Y => SharedReg797_out);

   SharedReg798_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg797_out,
                 Y => SharedReg798_out);

   SharedReg799_instance: Delay_34_DelayLength_56_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=56 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg798_out,
                 Y => SharedReg799_out);

   SharedReg800_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product710_3_impl_out,
                 Y => SharedReg800_out);

   SharedReg801_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg800_out,
                 Y => SharedReg801_out);

   SharedReg802_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg801_out,
                 Y => SharedReg802_out);

   SharedReg803_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg802_out,
                 Y => SharedReg803_out);

   SharedReg804_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg803_out,
                 Y => SharedReg804_out);

   SharedReg805_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg804_out,
                 Y => SharedReg805_out);

   SharedReg806_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg805_out,
                 Y => SharedReg806_out);

   SharedReg807_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg806_out,
                 Y => SharedReg807_out);

   SharedReg808_instance: Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=42 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg807_out,
                 Y => SharedReg808_out);

   SharedReg809_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product710_4_impl_out,
                 Y => SharedReg809_out);

   SharedReg810_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg809_out,
                 Y => SharedReg810_out);

   SharedReg811_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg810_out,
                 Y => SharedReg811_out);

   SharedReg812_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg811_out,
                 Y => SharedReg812_out);

   SharedReg813_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg812_out,
                 Y => SharedReg813_out);

   SharedReg814_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg813_out,
                 Y => SharedReg814_out);

   SharedReg815_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg814_out,
                 Y => SharedReg815_out);

   SharedReg816_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg815_out,
                 Y => SharedReg816_out);

   SharedReg817_instance: Delay_34_DelayLength_43_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=43 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg816_out,
                 Y => SharedReg817_out);

   SharedReg818_instance: Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=45 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg817_out,
                 Y => SharedReg818_out);

   SharedReg819_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product710_5_impl_out,
                 Y => SharedReg819_out);

   SharedReg820_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg819_out,
                 Y => SharedReg820_out);

   SharedReg821_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg820_out,
                 Y => SharedReg821_out);

   SharedReg822_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg821_out,
                 Y => SharedReg822_out);

   SharedReg823_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg822_out,
                 Y => SharedReg823_out);

   SharedReg824_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg823_out,
                 Y => SharedReg824_out);

   SharedReg825_instance: Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=44 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg824_out,
                 Y => SharedReg825_out);

   SharedReg826_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg825_out,
                 Y => SharedReg826_out);

   SharedReg827_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_0_impl_out,
                 Y => SharedReg827_out);

   SharedReg828_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg827_out,
                 Y => SharedReg828_out);

   SharedReg829_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg828_out,
                 Y => SharedReg829_out);

   SharedReg830_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg829_out,
                 Y => SharedReg830_out);

   SharedReg831_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg830_out,
                 Y => SharedReg831_out);

   SharedReg832_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg831_out,
                 Y => SharedReg832_out);

   SharedReg833_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg832_out,
                 Y => SharedReg833_out);

   SharedReg834_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg833_out,
                 Y => SharedReg834_out);

   SharedReg835_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_1_impl_out,
                 Y => SharedReg835_out);

   SharedReg836_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg835_out,
                 Y => SharedReg836_out);

   SharedReg837_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg836_out,
                 Y => SharedReg837_out);

   SharedReg838_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg837_out,
                 Y => SharedReg838_out);

   SharedReg839_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg838_out,
                 Y => SharedReg839_out);

   SharedReg840_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg839_out,
                 Y => SharedReg840_out);

   SharedReg841_instance: Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=40 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg840_out,
                 Y => SharedReg841_out);

   SharedReg842_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg841_out,
                 Y => SharedReg842_out);

   SharedReg843_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_2_impl_out,
                 Y => SharedReg843_out);

   SharedReg844_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg843_out,
                 Y => SharedReg844_out);

   SharedReg845_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg844_out,
                 Y => SharedReg845_out);

   SharedReg846_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg845_out,
                 Y => SharedReg846_out);

   SharedReg847_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg846_out,
                 Y => SharedReg847_out);

   SharedReg848_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg847_out,
                 Y => SharedReg848_out);

   SharedReg849_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg848_out,
                 Y => SharedReg849_out);

   SharedReg850_instance: Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=40 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg849_out,
                 Y => SharedReg850_out);

   SharedReg851_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg850_out,
                 Y => SharedReg851_out);

   SharedReg852_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_3_impl_out,
                 Y => SharedReg852_out);

   SharedReg853_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg852_out,
                 Y => SharedReg853_out);

   SharedReg854_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg853_out,
                 Y => SharedReg854_out);

   SharedReg855_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg854_out,
                 Y => SharedReg855_out);

   SharedReg856_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg855_out,
                 Y => SharedReg856_out);

   SharedReg857_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg856_out,
                 Y => SharedReg857_out);

   SharedReg858_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg857_out,
                 Y => SharedReg858_out);

   SharedReg859_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg858_out,
                 Y => SharedReg859_out);

   SharedReg860_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg859_out,
                 Y => SharedReg860_out);

   SharedReg861_instance: Delay_34_DelayLength_58_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=58 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg860_out,
                 Y => SharedReg861_out);

   SharedReg862_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_4_impl_out,
                 Y => SharedReg862_out);

   SharedReg863_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg862_out,
                 Y => SharedReg863_out);

   SharedReg864_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg863_out,
                 Y => SharedReg864_out);

   SharedReg865_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg864_out,
                 Y => SharedReg865_out);

   SharedReg866_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg865_out,
                 Y => SharedReg866_out);

   SharedReg867_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg866_out,
                 Y => SharedReg867_out);

   SharedReg868_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg867_out,
                 Y => SharedReg868_out);

   SharedReg869_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg868_out,
                 Y => SharedReg869_out);

   SharedReg870_instance: Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=31 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg869_out,
                 Y => SharedReg870_out);

   SharedReg871_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product810_5_impl_out,
                 Y => SharedReg871_out);

   SharedReg872_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg871_out,
                 Y => SharedReg872_out);

   SharedReg873_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg872_out,
                 Y => SharedReg873_out);

   SharedReg874_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg873_out,
                 Y => SharedReg874_out);

   SharedReg875_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg874_out,
                 Y => SharedReg875_out);

   SharedReg876_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg875_out,
                 Y => SharedReg876_out);

   SharedReg877_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg876_out,
                 Y => SharedReg877_out);

   SharedReg878_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg877_out,
                 Y => SharedReg878_out);

   SharedReg879_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product910_0_impl_out,
                 Y => SharedReg879_out);

   SharedReg880_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg879_out,
                 Y => SharedReg880_out);

   SharedReg881_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg880_out,
                 Y => SharedReg881_out);

   SharedReg882_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg881_out,
                 Y => SharedReg882_out);

   SharedReg883_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg882_out,
                 Y => SharedReg883_out);

   SharedReg884_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg883_out,
                 Y => SharedReg884_out);

   SharedReg885_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg884_out,
                 Y => SharedReg885_out);

   SharedReg886_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg885_out,
                 Y => SharedReg886_out);

   SharedReg887_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product910_1_impl_out,
                 Y => SharedReg887_out);

   SharedReg888_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg887_out,
                 Y => SharedReg888_out);

   SharedReg889_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg888_out,
                 Y => SharedReg889_out);

   SharedReg890_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg889_out,
                 Y => SharedReg890_out);

   SharedReg891_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg890_out,
                 Y => SharedReg891_out);

   SharedReg892_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg891_out,
                 Y => SharedReg892_out);

   SharedReg893_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product910_2_impl_out,
                 Y => SharedReg893_out);

   SharedReg894_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg893_out,
                 Y => SharedReg894_out);

   SharedReg895_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg894_out,
                 Y => SharedReg895_out);

   SharedReg896_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg895_out,
                 Y => SharedReg896_out);

   SharedReg897_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg896_out,
                 Y => SharedReg897_out);

   SharedReg898_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg897_out,
                 Y => SharedReg898_out);

   SharedReg899_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg898_out,
                 Y => SharedReg899_out);

   SharedReg900_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg899_out,
                 Y => SharedReg900_out);

   SharedReg901_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product910_3_impl_out,
                 Y => SharedReg901_out);

   SharedReg902_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg901_out,
                 Y => SharedReg902_out);

   SharedReg903_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg902_out,
                 Y => SharedReg903_out);

   SharedReg904_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg903_out,
                 Y => SharedReg904_out);

   SharedReg905_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg904_out,
                 Y => SharedReg905_out);

   SharedReg906_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg905_out,
                 Y => SharedReg906_out);

   SharedReg907_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product910_4_impl_out,
                 Y => SharedReg907_out);

   SharedReg908_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg907_out,
                 Y => SharedReg908_out);

   SharedReg909_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg908_out,
                 Y => SharedReg909_out);

   SharedReg910_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg909_out,
                 Y => SharedReg910_out);

   SharedReg911_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg910_out,
                 Y => SharedReg911_out);

   SharedReg912_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg911_out,
                 Y => SharedReg912_out);

   SharedReg913_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product910_5_impl_out,
                 Y => SharedReg913_out);

   SharedReg914_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg913_out,
                 Y => SharedReg914_out);

   SharedReg915_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg914_out,
                 Y => SharedReg915_out);

   SharedReg916_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg915_out,
                 Y => SharedReg916_out);

   SharedReg917_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg916_out,
                 Y => SharedReg917_out);

   SharedReg918_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg917_out,
                 Y => SharedReg918_out);

   SharedReg919_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg918_out,
                 Y => SharedReg919_out);

   SharedReg920_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg919_out,
                 Y => SharedReg920_out);

   SharedReg921_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg920_out,
                 Y => SharedReg921_out);

   SharedReg922_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg921_out,
                 Y => SharedReg922_out);

   SharedReg923_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg922_out,
                 Y => SharedReg923_out);

   SharedReg924_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_0_impl_out,
                 Y => SharedReg924_out);

   SharedReg925_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg924_out,
                 Y => SharedReg925_out);

   SharedReg926_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg925_out,
                 Y => SharedReg926_out);

   SharedReg927_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg926_out,
                 Y => SharedReg927_out);

   SharedReg928_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg927_out,
                 Y => SharedReg928_out);

   SharedReg929_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg928_out,
                 Y => SharedReg929_out);

   SharedReg930_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg929_out,
                 Y => SharedReg930_out);

   SharedReg931_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg930_out,
                 Y => SharedReg931_out);

   SharedReg932_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg931_out,
                 Y => SharedReg932_out);

   SharedReg933_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_1_impl_out,
                 Y => SharedReg933_out);

   SharedReg934_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg933_out,
                 Y => SharedReg934_out);

   SharedReg935_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg934_out,
                 Y => SharedReg935_out);

   SharedReg936_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg935_out,
                 Y => SharedReg936_out);

   SharedReg937_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg936_out,
                 Y => SharedReg937_out);

   SharedReg938_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg937_out,
                 Y => SharedReg938_out);

   SharedReg939_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg938_out,
                 Y => SharedReg939_out);

   SharedReg940_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg939_out,
                 Y => SharedReg940_out);

   SharedReg941_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg940_out,
                 Y => SharedReg941_out);

   SharedReg942_instance: Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=45 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg941_out,
                 Y => SharedReg942_out);

   SharedReg943_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_2_impl_out,
                 Y => SharedReg943_out);

   SharedReg944_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg943_out,
                 Y => SharedReg944_out);

   SharedReg945_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg944_out,
                 Y => SharedReg945_out);

   SharedReg946_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg945_out,
                 Y => SharedReg946_out);

   SharedReg947_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg946_out,
                 Y => SharedReg947_out);

   SharedReg948_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg947_out,
                 Y => SharedReg948_out);

   SharedReg949_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg948_out,
                 Y => SharedReg949_out);

   SharedReg950_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg949_out,
                 Y => SharedReg950_out);

   SharedReg951_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg950_out,
                 Y => SharedReg951_out);

   SharedReg952_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg951_out,
                 Y => SharedReg952_out);

   SharedReg953_instance: Delay_34_DelayLength_44_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=44 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg952_out,
                 Y => SharedReg953_out);

   SharedReg954_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg953_out,
                 Y => SharedReg954_out);

   SharedReg955_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg954_out,
                 Y => SharedReg955_out);

   SharedReg956_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_3_impl_out,
                 Y => SharedReg956_out);

   SharedReg957_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg956_out,
                 Y => SharedReg957_out);

   SharedReg958_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg957_out,
                 Y => SharedReg958_out);

   SharedReg959_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg958_out,
                 Y => SharedReg959_out);

   SharedReg960_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg959_out,
                 Y => SharedReg960_out);

   SharedReg961_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg960_out,
                 Y => SharedReg961_out);

   SharedReg962_instance: Delay_34_DelayLength_31_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=31 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg961_out,
                 Y => SharedReg962_out);

   SharedReg963_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg962_out,
                 Y => SharedReg963_out);

   SharedReg964_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg963_out,
                 Y => SharedReg964_out);

   SharedReg965_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_4_impl_out,
                 Y => SharedReg965_out);

   SharedReg966_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg965_out,
                 Y => SharedReg966_out);

   SharedReg967_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg966_out,
                 Y => SharedReg967_out);

   SharedReg968_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add30_5_impl_out,
                 Y => SharedReg968_out);

   SharedReg969_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg968_out,
                 Y => SharedReg969_out);

   SharedReg970_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg969_out,
                 Y => SharedReg970_out);

   SharedReg971_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg970_out,
                 Y => SharedReg971_out);

   SharedReg972_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg971_out,
                 Y => SharedReg972_out);

   SharedReg973_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg972_out,
                 Y => SharedReg973_out);

   SharedReg974_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg973_out,
                 Y => SharedReg974_out);

   SharedReg975_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg974_out,
                 Y => SharedReg975_out);

   SharedReg976_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg975_out,
                 Y => SharedReg976_out);

   SharedReg977_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add110_1_impl_out,
                 Y => SharedReg977_out);

   SharedReg978_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg977_out,
                 Y => SharedReg978_out);

   SharedReg979_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg978_out,
                 Y => SharedReg979_out);

   SharedReg980_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg979_out,
                 Y => SharedReg980_out);

   SharedReg981_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg980_out,
                 Y => SharedReg981_out);

   SharedReg982_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg981_out,
                 Y => SharedReg982_out);

   SharedReg983_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg982_out,
                 Y => SharedReg983_out);

   SharedReg984_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg983_out,
                 Y => SharedReg984_out);

   SharedReg985_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg984_out,
                 Y => SharedReg985_out);

   SharedReg986_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg985_out,
                 Y => SharedReg986_out);

   SharedReg987_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg986_out,
                 Y => SharedReg987_out);

   SharedReg988_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg987_out,
                 Y => SharedReg988_out);

   SharedReg989_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg988_out,
                 Y => SharedReg989_out);

   SharedReg990_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg989_out,
                 Y => SharedReg990_out);

   SharedReg991_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add110_2_impl_out,
                 Y => SharedReg991_out);

   SharedReg992_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg991_out,
                 Y => SharedReg992_out);

   SharedReg993_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg992_out,
                 Y => SharedReg993_out);

   SharedReg994_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg993_out,
                 Y => SharedReg994_out);

   SharedReg995_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg994_out,
                 Y => SharedReg995_out);

   SharedReg996_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg995_out,
                 Y => SharedReg996_out);

   SharedReg997_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg996_out,
                 Y => SharedReg997_out);

   SharedReg998_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg997_out,
                 Y => SharedReg998_out);

   SharedReg999_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg998_out,
                 Y => SharedReg999_out);

   SharedReg1000_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg999_out,
                 Y => SharedReg1000_out);

   SharedReg1001_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1000_out,
                 Y => SharedReg1001_out);

   SharedReg1002_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add110_3_impl_out,
                 Y => SharedReg1002_out);

   SharedReg1003_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1002_out,
                 Y => SharedReg1003_out);

   SharedReg1004_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1003_out,
                 Y => SharedReg1004_out);

   SharedReg1005_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1004_out,
                 Y => SharedReg1005_out);

   SharedReg1006_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1005_out,
                 Y => SharedReg1006_out);

   SharedReg1007_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1006_out,
                 Y => SharedReg1007_out);

   SharedReg1008_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1007_out,
                 Y => SharedReg1008_out);

   SharedReg1009_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1008_out,
                 Y => SharedReg1009_out);

   SharedReg1010_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1009_out,
                 Y => SharedReg1010_out);

   SharedReg1011_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add110_4_impl_out,
                 Y => SharedReg1011_out);

   SharedReg1012_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1011_out,
                 Y => SharedReg1012_out);

   SharedReg1013_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1012_out,
                 Y => SharedReg1013_out);

   SharedReg1014_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1013_out,
                 Y => SharedReg1014_out);

   SharedReg1015_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1014_out,
                 Y => SharedReg1015_out);

   SharedReg1016_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1015_out,
                 Y => SharedReg1016_out);

   SharedReg1017_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add101_2_impl_out,
                 Y => SharedReg1017_out);

   SharedReg1018_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1017_out,
                 Y => SharedReg1018_out);

   SharedReg1019_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1018_out,
                 Y => SharedReg1019_out);

   SharedReg1020_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1019_out,
                 Y => SharedReg1020_out);

   SharedReg1021_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1020_out,
                 Y => SharedReg1021_out);

   SharedReg1022_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1021_out,
                 Y => SharedReg1022_out);

   SharedReg1023_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1022_out,
                 Y => SharedReg1023_out);

   SharedReg1024_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1023_out,
                 Y => SharedReg1024_out);

   SharedReg1025_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1024_out,
                 Y => SharedReg1025_out);

   SharedReg1026_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1025_out,
                 Y => SharedReg1026_out);

   SharedReg1027_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1026_out,
                 Y => SharedReg1027_out);

   SharedReg1028_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add101_3_impl_out,
                 Y => SharedReg1028_out);

   SharedReg1029_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1028_out,
                 Y => SharedReg1029_out);

   SharedReg1030_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1029_out,
                 Y => SharedReg1030_out);

   SharedReg1031_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1030_out,
                 Y => SharedReg1031_out);

   SharedReg1032_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1031_out,
                 Y => SharedReg1032_out);

   SharedReg1033_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1032_out,
                 Y => SharedReg1033_out);

   SharedReg1034_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1033_out,
                 Y => SharedReg1034_out);

   SharedReg1035_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1034_out,
                 Y => SharedReg1035_out);

   SharedReg1036_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1035_out,
                 Y => SharedReg1036_out);

   SharedReg1037_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1036_out,
                 Y => SharedReg1037_out);

   SharedReg1038_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1037_out,
                 Y => SharedReg1038_out);

   SharedReg1039_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1038_out,
                 Y => SharedReg1039_out);

   SharedReg1040_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1039_out,
                 Y => SharedReg1040_out);

   SharedReg1041_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1040_out,
                 Y => SharedReg1041_out);

   SharedReg1042_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1041_out,
                 Y => SharedReg1042_out);

   SharedReg1043_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1042_out,
                 Y => SharedReg1043_out);

   SharedReg1044_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add101_5_impl_out,
                 Y => SharedReg1044_out);

   SharedReg1045_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1044_out,
                 Y => SharedReg1045_out);

   SharedReg1046_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1045_out,
                 Y => SharedReg1046_out);

   SharedReg1047_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1046_out,
                 Y => SharedReg1047_out);

   SharedReg1048_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1047_out,
                 Y => SharedReg1048_out);

   SharedReg1049_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1048_out,
                 Y => SharedReg1049_out);

   SharedReg1050_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1049_out,
                 Y => SharedReg1050_out);

   SharedReg1051_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1050_out,
                 Y => SharedReg1051_out);

   SharedReg1052_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1051_out,
                 Y => SharedReg1052_out);

   SharedReg1053_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1052_out,
                 Y => SharedReg1053_out);

   SharedReg1054_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1053_out,
                 Y => SharedReg1054_out);

   SharedReg1055_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1054_out,
                 Y => SharedReg1055_out);

   SharedReg1056_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1055_out,
                 Y => SharedReg1056_out);

   SharedReg1057_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1056_out,
                 Y => SharedReg1057_out);

   SharedReg1058_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1057_out,
                 Y => SharedReg1058_out);

   SharedReg1059_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add111_1_impl_out,
                 Y => SharedReg1059_out);

   SharedReg1060_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1059_out,
                 Y => SharedReg1060_out);

   SharedReg1061_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1060_out,
                 Y => SharedReg1061_out);

   SharedReg1062_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1061_out,
                 Y => SharedReg1062_out);

   SharedReg1063_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1062_out,
                 Y => SharedReg1063_out);

   SharedReg1064_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1063_out,
                 Y => SharedReg1064_out);

   SharedReg1065_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1064_out,
                 Y => SharedReg1065_out);

   SharedReg1066_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1065_out,
                 Y => SharedReg1066_out);

   SharedReg1067_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1066_out,
                 Y => SharedReg1067_out);

   SharedReg1068_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1067_out,
                 Y => SharedReg1068_out);

   SharedReg1069_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1068_out,
                 Y => SharedReg1069_out);

   SharedReg1070_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add111_4_impl_out,
                 Y => SharedReg1070_out);

   SharedReg1071_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1070_out,
                 Y => SharedReg1071_out);

   SharedReg1072_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1071_out,
                 Y => SharedReg1072_out);

   SharedReg1073_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1072_out,
                 Y => SharedReg1073_out);

   SharedReg1074_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1073_out,
                 Y => SharedReg1074_out);

   SharedReg1075_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1074_out,
                 Y => SharedReg1075_out);

   SharedReg1076_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1075_out,
                 Y => SharedReg1076_out);

   SharedReg1077_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1076_out,
                 Y => SharedReg1077_out);

   SharedReg1078_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1077_out,
                 Y => SharedReg1078_out);

   SharedReg1079_instance: Delay_34_DelayLength_40_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=40 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1078_out,
                 Y => SharedReg1079_out);

   SharedReg1080_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1079_out,
                 Y => SharedReg1080_out);

   SharedReg1081_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1080_out,
                 Y => SharedReg1081_out);

   SharedReg1082_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add141_0_impl_out,
                 Y => SharedReg1082_out);

   SharedReg1083_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1082_out,
                 Y => SharedReg1083_out);

   SharedReg1084_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1083_out,
                 Y => SharedReg1084_out);

   SharedReg1085_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1084_out,
                 Y => SharedReg1085_out);

   SharedReg1086_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1085_out,
                 Y => SharedReg1086_out);

   SharedReg1087_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1086_out,
                 Y => SharedReg1087_out);

   SharedReg1088_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1087_out,
                 Y => SharedReg1088_out);

   SharedReg1089_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1088_out,
                 Y => SharedReg1089_out);

   SharedReg1090_instance: Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=45 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1089_out,
                 Y => SharedReg1090_out);

   SharedReg1091_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add141_2_impl_out,
                 Y => SharedReg1091_out);

   SharedReg1092_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1091_out,
                 Y => SharedReg1092_out);

   SharedReg1093_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1092_out,
                 Y => SharedReg1093_out);

   SharedReg1094_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add141_3_impl_out,
                 Y => SharedReg1094_out);

   SharedReg1095_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1094_out,
                 Y => SharedReg1095_out);

   SharedReg1096_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1095_out,
                 Y => SharedReg1096_out);

   SharedReg1097_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1096_out,
                 Y => SharedReg1097_out);

   SharedReg1098_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1097_out,
                 Y => SharedReg1098_out);

   SharedReg1099_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1098_out,
                 Y => SharedReg1099_out);

   SharedReg1100_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1099_out,
                 Y => SharedReg1100_out);

   SharedReg1101_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1100_out,
                 Y => SharedReg1101_out);

   SharedReg1102_instance: Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=50 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1101_out,
                 Y => SharedReg1102_out);

   SharedReg1103_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1102_out,
                 Y => SharedReg1103_out);

   SharedReg1104_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add141_5_impl_out,
                 Y => SharedReg1104_out);

   SharedReg1105_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1104_out,
                 Y => SharedReg1105_out);

   SharedReg1106_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1105_out,
                 Y => SharedReg1106_out);

   SharedReg1107_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1106_out,
                 Y => SharedReg1107_out);

   SharedReg1108_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1107_out,
                 Y => SharedReg1108_out);

   SharedReg1109_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1108_out,
                 Y => SharedReg1109_out);

   SharedReg1110_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1109_out,
                 Y => SharedReg1110_out);

   SharedReg1111_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1110_out,
                 Y => SharedReg1111_out);

   SharedReg1112_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1111_out,
                 Y => SharedReg1112_out);

   SharedReg1113_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1112_out,
                 Y => SharedReg1113_out);

   SharedReg1114_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1113_out,
                 Y => SharedReg1114_out);

   SharedReg1115_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add151_5_impl_out,
                 Y => SharedReg1115_out);

   SharedReg1116_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1115_out,
                 Y => SharedReg1116_out);

   SharedReg1117_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1116_out,
                 Y => SharedReg1117_out);

   SharedReg1118_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1117_out,
                 Y => SharedReg1118_out);

   SharedReg1119_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1118_out,
                 Y => SharedReg1119_out);

   SharedReg1120_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1119_out,
                 Y => SharedReg1120_out);

   SharedReg1121_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1120_out,
                 Y => SharedReg1121_out);

   SharedReg1122_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1121_out,
                 Y => SharedReg1122_out);

   SharedReg1123_instance: Delay_34_DelayLength_50_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=50 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1122_out,
                 Y => SharedReg1123_out);

   SharedReg1124_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1123_out,
                 Y => SharedReg1124_out);

   SharedReg1125_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1124_out,
                 Y => SharedReg1125_out);

   SharedReg1126_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1125_out,
                 Y => SharedReg1126_out);

   SharedReg1127_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add21_3_impl_out,
                 Y => SharedReg1127_out);

   SharedReg1128_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1127_out,
                 Y => SharedReg1128_out);

   SharedReg1129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1128_out,
                 Y => SharedReg1129_out);

   SharedReg1130_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1129_out,
                 Y => SharedReg1130_out);

   SharedReg1131_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1130_out,
                 Y => SharedReg1131_out);

   SharedReg1132_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1131_out,
                 Y => SharedReg1132_out);

   SharedReg1133_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1132_out,
                 Y => SharedReg1133_out);

   SharedReg1134_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1133_out,
                 Y => SharedReg1134_out);

   SharedReg1135_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1134_out,
                 Y => SharedReg1135_out);

   SharedReg1136_instance: Delay_34_DelayLength_45_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=45 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1135_out,
                 Y => SharedReg1136_out);

   SharedReg1137_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add23_0_impl_out,
                 Y => SharedReg1137_out);

   SharedReg1138_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1137_out,
                 Y => SharedReg1138_out);

   SharedReg1139_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1138_out,
                 Y => SharedReg1139_out);

   SharedReg1140_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1139_out,
                 Y => SharedReg1140_out);

   SharedReg1141_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1140_out,
                 Y => SharedReg1141_out);

   SharedReg1142_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1141_out,
                 Y => SharedReg1142_out);

   SharedReg1143_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1142_out,
                 Y => SharedReg1143_out);

   SharedReg1144_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1143_out,
                 Y => SharedReg1144_out);

   SharedReg1145_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1144_out,
                 Y => SharedReg1145_out);

   SharedReg1146_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1145_out,
                 Y => SharedReg1146_out);

   SharedReg1147_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1146_out,
                 Y => SharedReg1147_out);

   SharedReg1148_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product312_0_impl_out,
                 Y => SharedReg1148_out);

   SharedReg1149_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1148_out,
                 Y => SharedReg1149_out);

   SharedReg1150_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1149_out,
                 Y => SharedReg1150_out);

   SharedReg1151_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1150_out,
                 Y => SharedReg1151_out);

   SharedReg1152_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1151_out,
                 Y => SharedReg1152_out);

   SharedReg1153_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product312_1_impl_out,
                 Y => SharedReg1153_out);

   SharedReg1154_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1153_out,
                 Y => SharedReg1154_out);

   SharedReg1155_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1154_out,
                 Y => SharedReg1155_out);

   SharedReg1156_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1155_out,
                 Y => SharedReg1156_out);

   SharedReg1157_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1156_out,
                 Y => SharedReg1157_out);

   SharedReg1158_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1157_out,
                 Y => SharedReg1158_out);

   SharedReg1159_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1158_out,
                 Y => SharedReg1159_out);

   SharedReg1160_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product312_2_impl_out,
                 Y => SharedReg1160_out);

   SharedReg1161_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1160_out,
                 Y => SharedReg1161_out);

   SharedReg1162_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1161_out,
                 Y => SharedReg1162_out);

   SharedReg1163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1162_out,
                 Y => SharedReg1163_out);

   SharedReg1164_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1163_out,
                 Y => SharedReg1164_out);

   SharedReg1165_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1164_out,
                 Y => SharedReg1165_out);

   SharedReg1166_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1165_out,
                 Y => SharedReg1166_out);

   SharedReg1167_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product312_3_impl_out,
                 Y => SharedReg1167_out);

   SharedReg1168_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1167_out,
                 Y => SharedReg1168_out);

   SharedReg1169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1168_out,
                 Y => SharedReg1169_out);

   SharedReg1170_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1169_out,
                 Y => SharedReg1170_out);

   SharedReg1171_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1170_out,
                 Y => SharedReg1171_out);

   SharedReg1172_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1171_out,
                 Y => SharedReg1172_out);

   SharedReg1173_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1172_out,
                 Y => SharedReg1173_out);

   SharedReg1174_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product312_4_impl_out,
                 Y => SharedReg1174_out);

   SharedReg1175_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1174_out,
                 Y => SharedReg1175_out);

   SharedReg1176_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1175_out,
                 Y => SharedReg1176_out);

   SharedReg1177_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1176_out,
                 Y => SharedReg1177_out);

   SharedReg1178_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1177_out,
                 Y => SharedReg1178_out);

   SharedReg1179_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1178_out,
                 Y => SharedReg1179_out);

   SharedReg1180_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1179_out,
                 Y => SharedReg1180_out);

   SharedReg1181_instance: Delay_34_DelayLength_49_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=49 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1180_out,
                 Y => SharedReg1181_out);

   SharedReg1182_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1181_out,
                 Y => SharedReg1182_out);

   SharedReg1183_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product312_5_impl_out,
                 Y => SharedReg1183_out);

   SharedReg1184_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1183_out,
                 Y => SharedReg1184_out);

   SharedReg1185_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1184_out,
                 Y => SharedReg1185_out);

   SharedReg1186_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1185_out,
                 Y => SharedReg1186_out);

   SharedReg1187_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1186_out,
                 Y => SharedReg1187_out);

   SharedReg1188_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1187_out,
                 Y => SharedReg1188_out);

   SharedReg1189_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1188_out,
                 Y => SharedReg1189_out);

   SharedReg1190_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1189_out,
                 Y => SharedReg1190_out);

   SharedReg1191_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product54_4_impl_out,
                 Y => SharedReg1191_out);

   SharedReg1192_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1191_out,
                 Y => SharedReg1192_out);

   SharedReg1193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1192_out,
                 Y => SharedReg1193_out);

   SharedReg1194_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1193_out,
                 Y => SharedReg1194_out);

   SharedReg1195_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1194_out,
                 Y => SharedReg1195_out);

   SharedReg1196_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1195_out,
                 Y => SharedReg1196_out);

   SharedReg1197_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1196_out,
                 Y => SharedReg1197_out);

   SharedReg1198_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1197_out,
                 Y => SharedReg1198_out);

   SharedReg1199_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1198_out,
                 Y => SharedReg1199_out);

   SharedReg1200_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product54_5_impl_out,
                 Y => SharedReg1200_out);

   SharedReg1201_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1200_out,
                 Y => SharedReg1201_out);

   SharedReg1202_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1201_out,
                 Y => SharedReg1202_out);

   SharedReg1203_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1202_out,
                 Y => SharedReg1203_out);

   SharedReg1204_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1203_out,
                 Y => SharedReg1204_out);

   SharedReg1205_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1204_out,
                 Y => SharedReg1205_out);

   SharedReg1206_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1205_out,
                 Y => SharedReg1206_out);

   SharedReg1207_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product62_5_impl_out,
                 Y => SharedReg1207_out);

   SharedReg1208_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1207_out,
                 Y => SharedReg1208_out);

   SharedReg1209_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1208_out,
                 Y => SharedReg1209_out);

   SharedReg1210_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1209_out,
                 Y => SharedReg1210_out);

   SharedReg1211_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1210_out,
                 Y => SharedReg1211_out);

   SharedReg1212_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_0_impl_out,
                 Y => SharedReg1212_out);

   SharedReg1213_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1212_out,
                 Y => SharedReg1213_out);

   SharedReg1214_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1213_out,
                 Y => SharedReg1214_out);

   SharedReg1215_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1214_out,
                 Y => SharedReg1215_out);

   SharedReg1216_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1215_out,
                 Y => SharedReg1216_out);

   SharedReg1217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1216_out,
                 Y => SharedReg1217_out);

   SharedReg1218_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_1_impl_out,
                 Y => SharedReg1218_out);

   SharedReg1219_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1218_out,
                 Y => SharedReg1219_out);

   SharedReg1220_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1219_out,
                 Y => SharedReg1220_out);

   SharedReg1221_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1220_out,
                 Y => SharedReg1221_out);

   SharedReg1222_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1221_out,
                 Y => SharedReg1222_out);

   SharedReg1223_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1222_out,
                 Y => SharedReg1223_out);

   SharedReg1224_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_2_impl_out,
                 Y => SharedReg1224_out);

   SharedReg1225_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1224_out,
                 Y => SharedReg1225_out);

   SharedReg1226_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1225_out,
                 Y => SharedReg1226_out);

   SharedReg1227_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1226_out,
                 Y => SharedReg1227_out);

   SharedReg1228_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1227_out,
                 Y => SharedReg1228_out);

   SharedReg1229_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1228_out,
                 Y => SharedReg1229_out);

   SharedReg1230_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_3_impl_out,
                 Y => SharedReg1230_out);

   SharedReg1231_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1230_out,
                 Y => SharedReg1231_out);

   SharedReg1232_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1231_out,
                 Y => SharedReg1232_out);

   SharedReg1233_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1232_out,
                 Y => SharedReg1233_out);

   SharedReg1234_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1233_out,
                 Y => SharedReg1234_out);

   SharedReg1235_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1234_out,
                 Y => SharedReg1235_out);

   SharedReg1236_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_4_impl_out,
                 Y => SharedReg1236_out);

   SharedReg1237_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1236_out,
                 Y => SharedReg1237_out);

   SharedReg1238_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1237_out,
                 Y => SharedReg1238_out);

   SharedReg1239_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1238_out,
                 Y => SharedReg1239_out);

   SharedReg1240_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1239_out,
                 Y => SharedReg1240_out);

   SharedReg1241_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1240_out,
                 Y => SharedReg1241_out);

   SharedReg1242_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Subtract12_5_impl_out,
                 Y => SharedReg1242_out);

   SharedReg1243_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1242_out,
                 Y => SharedReg1243_out);

   SharedReg1244_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1243_out,
                 Y => SharedReg1244_out);

   SharedReg1245_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1244_out,
                 Y => SharedReg1245_out);

   SharedReg1246_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1245_out,
                 Y => SharedReg1246_out);

   SharedReg1247_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1246_out,
                 Y => SharedReg1247_out);

   SharedReg1248_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Add10_5_impl_out,
                 Y => SharedReg1248_out);

   SharedReg1249_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1248_out,
                 Y => SharedReg1249_out);

   SharedReg1250_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1249_out,
                 Y => SharedReg1250_out);

   SharedReg1251_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1250_out,
                 Y => SharedReg1251_out);

   SharedReg1252_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1251_out,
                 Y => SharedReg1252_out);

   SharedReg1253_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1252_out,
                 Y => SharedReg1253_out);

   SharedReg1254_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1253_out,
                 Y => SharedReg1254_out);

   SharedReg1255_instance: Delay_34_DelayLength_103_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=103 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_0_impl_out,
                 Y => SharedReg1255_out);

   SharedReg1256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Divide_0_impl_out,
                 Y => SharedReg1256_out);

   SharedReg1257_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product213_5_impl_out,
                 Y => SharedReg1257_out);

   SharedReg1258_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1257_out,
                 Y => SharedReg1258_out);

   SharedReg1259_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1258_out,
                 Y => SharedReg1259_out);

   SharedReg1260_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1259_out,
                 Y => SharedReg1260_out);

   SharedReg1261_instance: Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=42 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1260_out,
                 Y => SharedReg1261_out);

   SharedReg1262_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1261_out,
                 Y => SharedReg1262_out);

   SharedReg1263_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_0_impl_out,
                 Y => SharedReg1263_out);

   SharedReg1264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1263_out,
                 Y => SharedReg1264_out);

   SharedReg1265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1264_out,
                 Y => SharedReg1265_out);

   SharedReg1266_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1265_out,
                 Y => SharedReg1266_out);

   SharedReg1267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1266_out,
                 Y => SharedReg1267_out);

   SharedReg1268_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1267_out,
                 Y => SharedReg1268_out);

   SharedReg1269_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1268_out,
                 Y => SharedReg1269_out);

   SharedReg1270_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1269_out,
                 Y => SharedReg1270_out);

   SharedReg1271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1270_out,
                 Y => SharedReg1271_out);

   SharedReg1272_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1271_out,
                 Y => SharedReg1272_out);

   SharedReg1273_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1272_out,
                 Y => SharedReg1273_out);

   SharedReg1274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1273_out,
                 Y => SharedReg1274_out);

   SharedReg1275_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1274_out,
                 Y => SharedReg1275_out);

   SharedReg1276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1275_out,
                 Y => SharedReg1276_out);

   SharedReg1277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1276_out,
                 Y => SharedReg1277_out);

   SharedReg1278_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1277_out,
                 Y => SharedReg1278_out);

   SharedReg1279_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1278_out,
                 Y => SharedReg1279_out);

   SharedReg1280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1279_out,
                 Y => SharedReg1280_out);

   SharedReg1281_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1280_out,
                 Y => SharedReg1281_out);

   SharedReg1282_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1281_out,
                 Y => SharedReg1282_out);

   SharedReg1283_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1282_out,
                 Y => SharedReg1283_out);

   SharedReg1284_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1283_out,
                 Y => SharedReg1284_out);

   SharedReg1285_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1284_out,
                 Y => SharedReg1285_out);

   SharedReg1286_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1285_out,
                 Y => SharedReg1286_out);

   SharedReg1287_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1286_out,
                 Y => SharedReg1287_out);

   SharedReg1288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1287_out,
                 Y => SharedReg1288_out);

   SharedReg1289_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1288_out,
                 Y => SharedReg1289_out);

   SharedReg1290_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1289_out,
                 Y => SharedReg1290_out);

   SharedReg1291_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1290_out,
                 Y => SharedReg1291_out);

   SharedReg1292_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1291_out,
                 Y => SharedReg1292_out);

   SharedReg1293_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1292_out,
                 Y => SharedReg1293_out);

   SharedReg1294_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1293_out,
                 Y => SharedReg1294_out);

   SharedReg1295_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1294_out,
                 Y => SharedReg1295_out);

   SharedReg1296_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1295_out,
                 Y => SharedReg1296_out);

   SharedReg1297_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1296_out,
                 Y => SharedReg1297_out);

   SharedReg1298_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1297_out,
                 Y => SharedReg1298_out);

   SharedReg1299_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1298_out,
                 Y => SharedReg1299_out);

   SharedReg1300_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1299_out,
                 Y => SharedReg1300_out);

   SharedReg1301_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1300_out,
                 Y => SharedReg1301_out);

   SharedReg1302_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1301_out,
                 Y => SharedReg1302_out);

   SharedReg1303_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1302_out,
                 Y => SharedReg1303_out);

   SharedReg1304_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1303_out,
                 Y => SharedReg1304_out);

   SharedReg1305_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1304_out,
                 Y => SharedReg1305_out);

   SharedReg1306_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1305_out,
                 Y => SharedReg1306_out);

   SharedReg1307_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1306_out,
                 Y => SharedReg1307_out);

   SharedReg1308_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1307_out,
                 Y => SharedReg1308_out);

   SharedReg1309_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1308_out,
                 Y => SharedReg1309_out);

   SharedReg1310_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1309_out,
                 Y => SharedReg1310_out);

   SharedReg1311_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1310_out,
                 Y => SharedReg1311_out);

   SharedReg1312_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1311_out,
                 Y => SharedReg1312_out);

   SharedReg1313_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1312_out,
                 Y => SharedReg1313_out);

   SharedReg1314_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1313_out,
                 Y => SharedReg1314_out);

   SharedReg1315_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1314_out,
                 Y => SharedReg1315_out);

   SharedReg1316_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1315_out,
                 Y => SharedReg1316_out);

   SharedReg1317_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1316_out,
                 Y => SharedReg1317_out);
end architecture;

