--------------------------------------------------------------------------------
--                         ModuloCounter_59_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity ModuloCounter_59_component is
   port ( clk, rst : in std_logic;
          Counter_out : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of ModuloCounter_59_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk,rst)
	 variable count : std_logic_vector(5 downto 0) := (others => '0');
begin
	 if rst = '1' then
	 	 count := (others => '0');
	 elsif clk'event and clk = '1' then
	 	 if count = 58 then
	 	 	 count := (others => '0');
	 	 else
	 	 	 count := count+1;
	 	 end if;
	 end if;
	 Counter_out <= count;
end process;
end architecture;

--------------------------------------------------------------------------------
--                          InputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(31 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of InputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal expInfty : std_logic := '0';
signal fracZero : std_logic := '0';
signal reprSubNormal : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal infinity : std_logic := '0';
signal zero : std_logic := '0';
signal NaN : std_logic := '0';
signal exnR : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_31_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_31_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_31_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111001111110000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_28_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_28_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_28_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111001111000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n352_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n352_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n352_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111011101100000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n432_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n432_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n432_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111011110110000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n500_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n500_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n500_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111011111110100000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n532_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n532_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n532_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111100000001010000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n129_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n129_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n129_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111011000000010000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_158_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_158_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_158_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111011000111100000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_526_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_526_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_526_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111100000000111000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_964_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_964_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_964_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111100011100010000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n529_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n529_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n529_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111100000001000100000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n464_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n464_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n464_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111011111010000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_29_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_29_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_29_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111001111010000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n336_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n336_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n336_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111011101010000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_3136_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_3136_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_3136_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111101010001000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_3648_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_3648_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_3648_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111101011001000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_4110_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_4110_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_4110_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111101100000000111000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_4478_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_4478_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_4478_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111101100010111111000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_4737_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_4737_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_4737_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111101100101000000100000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_4868_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_4868_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_4868_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111101100110000010000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_22_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_22_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_22_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111001101100000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_1472_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_1472_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_1472_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111100101110000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_2008_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_2008_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_2008_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111100111110110000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_2576_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_2576_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_2576_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111101001000010000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                 Constant_float_8_23_8_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_8_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_8_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0100111001000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n17_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n17_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n17_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111001100010000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n59_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n59_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n59_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111010011011000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n116_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n116_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n116_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111010111010000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n188_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n188_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n188_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111011001111000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                Constant_float_8_23_n268_div_65536_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Patrick Sittel
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Constant_float_8_23_n268_div_65536_component is
   port ( clk, rst : in std_logic;
          Y : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of Constant_float_8_23_n268_div_65536_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
---------------------  addFullComment for a large comment  ---------------------
   -- addComment for small left-aligned comment
    Y <= "0110111011100001100000000000000000";
end architecture;

--------------------------------------------------------------------------------
--          IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid6324599
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid6324599 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          Y : in std_logic_vector(23 downto 0);
          R : out std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid6324599 is
signal XX_m6324600 : std_logic_vector(23 downto 0) := (others => '0');
signal YY_m6324600 : std_logic_vector(23 downto 0) := (others => '0');
signal XX : unsigned(-1+24 downto 0) := (others => '0');
signal YY : unsigned(-1+24 downto 0) := (others => '0');
signal RR : unsigned(-1+48 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   XX_m6324600 <= X ;
   YY_m6324600 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(47 downto 0));
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_33_f500_uid6324603
--                   (IntAdderClassical_33_f500_uid6324605)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f500_uid6324603 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(32 downto 0);
          Y : in std_logic_vector(32 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f500_uid6324603 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--         FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid6324599 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             Y : in std_logic_vector(23 downto 0);
             R : out std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f500_uid6324603 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(32 downto 0);
             Y : in std_logic_vector(32 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 : std_logic := '0';
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal expY : std_logic_vector(7 downto 0) := (others => '0');
signal expSumPreSub, expSumPreSub_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal bias, bias_d1 : std_logic_vector(9 downto 0) := (others => '0');
signal expSum : std_logic_vector(9 downto 0) := (others => '0');
signal sigX : std_logic_vector(23 downto 0) := (others => '0');
signal sigY : std_logic_vector(23 downto 0) := (others => '0');
signal sigProd, sigProd_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal excSel : std_logic_vector(3 downto 0) := (others => '0');
signal exc, exc_d1, exc_d2 : std_logic_vector(1 downto 0) := (others => '0');
signal norm : std_logic := '0';
signal expPostNorm : std_logic_vector(9 downto 0) := (others => '0');
signal sigProdExt, sigProdExt_d1 : std_logic_vector(47 downto 0) := (others => '0');
signal expSig, expSig_d1 : std_logic_vector(32 downto 0) := (others => '0');
signal sticky, sticky_d1 : std_logic := '0';
signal guard, guard_d1 : std_logic := '0';
signal round : std_logic := '0';
signal expSigPostRound : std_logic_vector(32 downto 0) := (others => '0');
signal excPostNorm : std_logic_vector(1 downto 0) := (others => '0');
signal finalExc : std_logic_vector(1 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
            guard_d1 <=  guard;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   ----------------Synchro barrier, entering cycle 1----------------
   expSum <= expSumPreSub_d1 - bias_d1;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F500_uid6324599  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd_d1(47);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(46 downto 0) & "0" when norm='1' else
                         sigProd_d1(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   ----------------Synchro barrier, entering cycle 2----------------
   round <= sticky_d1 and ( (guard_d1 and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
      RoundingAdder: IntAdder_33_f500_uid6324603  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_55_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_55_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iS_47 : in std_logic_vector(33 downto 0);
          iS_48 : in std_logic_vector(33 downto 0);
          iS_49 : in std_logic_vector(33 downto 0);
          iS_50 : in std_logic_vector(33 downto 0);
          iS_51 : in std_logic_vector(33 downto 0);
          iS_52 : in std_logic_vector(33 downto 0);
          iS_53 : in std_logic_vector(33 downto 0);
          iS_54 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_55_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
         iS_47 when "101111",
         iS_48 when "110000",
         iS_49 when "110001",
         iS_50 when "110010",
         iS_51 when "110011",
         iS_52 when "110100",
         iS_53 when "110101",
         iS_54 when "110110",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      Y <= s0;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_41_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_41_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_41_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_19_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_19_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(4 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_19_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "00000",
         iS_1 when "00001",
         iS_2 when "00010",
         iS_3 when "00011",
         iS_4 when "00100",
         iS_5 when "00101",
         iS_6 when "00110",
         iS_7 when "00111",
         iS_8 when "01000",
         iS_9 when "01001",
         iS_10 when "01010",
         iS_11 when "01011",
         iS_12 when "01100",
         iS_13 when "01101",
         iS_14 when "01110",
         iS_15 when "01111",
         iS_16 when "10000",
         iS_17 when "10001",
         iS_18 when "10010",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_5_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_5_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(2 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_5_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000",
         iS_1 when "001",
         iS_2 when "010",
         iS_3 when "011",
         iS_4 when "100",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                     FPAdd_8_23_uid6324686_RightShifter
--                (RightShifter_24_by_max_26_F250_uid6324688)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid6324686_RightShifter is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(23 downto 0);
          S : in std_logic_vector(4 downto 0);
          R : out std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid6324686_RightShifter is
signal level0 : std_logic_vector(23 downto 0) := (others => '0');
signal ps : std_logic_vector(4 downto 0) := (others => '0');
signal level1 : std_logic_vector(24 downto 0) := (others => '0');
signal level2 : std_logic_vector(26 downto 0) := (others => '0');
signal level3 : std_logic_vector(30 downto 0) := (others => '0');
signal level4 : std_logic_vector(38 downto 0) := (others => '0');
signal level5 : std_logic_vector(54 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(54 downto 5);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_27_f250_uid6324691
--                  (IntAdderAlternative_27_f250_uid6324695)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_f250_uid6324691 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(26 downto 0);
          Y : in std_logic_vector(26 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_f250_uid6324691 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--              LZCShifter_28_to_28_counting_32_F250_uid6324698
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_28_to_28_counting_32_F250_uid6324698 is
   port ( clk, rst : in std_logic;
          I : in std_logic_vector(27 downto 0);
          Count : out std_logic_vector(4 downto 0);
          O : out std_logic_vector(27 downto 0)   );
end entity;

architecture arch of LZCShifter_28_to_28_counting_32_F250_uid6324698 is
signal level5 : std_logic_vector(27 downto 0) := (others => '0');
signal count4, count4_d1 : std_logic := '0';
signal level4, level4_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal count3, count3_d1 : std_logic := '0';
signal level3 : std_logic_vector(27 downto 0) := (others => '0');
signal count2 : std_logic := '0';
signal level2 : std_logic_vector(27 downto 0) := (others => '0');
signal count1 : std_logic := '0';
signal level1 : std_logic_vector(27 downto 0) := (others => '0');
signal count0 : std_logic := '0';
signal level0 : std_logic_vector(27 downto 0) := (others => '0');
signal sCount : std_logic_vector(4 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
         end if;
      end process;
   level5 <= I ;
   count4<= '1' when level5(27 downto 12) = (27 downto 12=>'0') else '0';
   level4<= level5(27 downto 0) when count4='0' else level5(11 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(27 downto 20) = (27 downto 20=>'0') else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level4_d1(27 downto 0) when count3_d1='0' else level4_d1(19 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(27 downto 24) = (27 downto 24=>'0') else '0';
   level2<= level3(27 downto 0) when count2='0' else level3(23 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(27 downto 26) = (27 downto 26=>'0') else '0';
   level1<= level2(27 downto 0) when count1='0' else level2(25 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0<= level1(27 downto 0) when count0='0' else level1(26 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count4_d1 & count3_d1 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_34_f250_uid6324701
--                   (IntAdderClassical_34_f250_uid6324703)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_f250_uid6324701 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : in std_logic_vector(33 downto 0);
          Cin : in std_logic;
          R : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_f250_uid6324701 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                           FPAdd_8_23_uid6324686
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdd_8_23_uid6324686 is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPAdd_8_23_uid6324686 is
   component FPAdd_8_23_uid6324686_RightShifter is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(23 downto 0);
             S : in std_logic_vector(4 downto 0);
             R : out std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_27_f250_uid6324691 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(26 downto 0);
             Y : in std_logic_vector(26 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(26 downto 0)   );
   end component;

   component LZCShifter_28_to_28_counting_32_F250_uid6324698 is
      port ( clk, rst : in std_logic;
             I : in std_logic_vector(27 downto 0);
             Count : out std_logic_vector(4 downto 0);
             O : out std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_f250_uid6324701 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : in std_logic_vector(33 downto 0);
             Cin : in std_logic;
             R : out std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX : std_logic_vector(32 downto 0) := (others => '0');
signal excExpFracY : std_logic_vector(32 downto 0) := (others => '0');
signal eXmeY : std_logic_vector(8 downto 0) := (others => '0');
signal eYmeX : std_logic_vector(8 downto 0) := (others => '0');
signal swap : std_logic := '0';
signal newX, newX_d1 : std_logic_vector(33 downto 0) := (others => '0');
signal newY : std_logic_vector(33 downto 0) := (others => '0');
signal expX, expX_d1 : std_logic_vector(7 downto 0) := (others => '0');
signal excX : std_logic_vector(1 downto 0) := (others => '0');
signal excY : std_logic_vector(1 downto 0) := (others => '0');
signal signX : std_logic := '0';
signal signY : std_logic := '0';
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3 : std_logic := '0';
signal sXsYExnXY : std_logic_vector(5 downto 0) := (others => '0');
signal sdExnXY : std_logic_vector(3 downto 0) := (others => '0');
signal fracY : std_logic_vector(23 downto 0) := (others => '0');
signal excRt, excRt_d1, excRt_d2, excRt_d3 : std_logic_vector(1 downto 0) := (others => '0');
signal signR, signR_d1, signR_d2, signR_d3 : std_logic := '0';
signal expDiff : std_logic_vector(8 downto 0) := (others => '0');
signal shiftedOut : std_logic := '0';
signal shiftVal : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFracY, shiftedFracY_d1 : std_logic_vector(49 downto 0) := (others => '0');
signal sticky : std_logic := '0';
signal fracYfar : std_logic_vector(26 downto 0) := (others => '0');
signal EffSubVector : std_logic_vector(26 downto 0) := (others => '0');
signal fracYfarXorOp : std_logic_vector(26 downto 0) := (others => '0');
signal fracXfar : std_logic_vector(26 downto 0) := (others => '0');
signal cInAddFar : std_logic := '0';
signal fracAddResult : std_logic_vector(26 downto 0) := (others => '0');
signal fracGRS : std_logic_vector(27 downto 0) := (others => '0');
signal extendedExpInc, extendedExpInc_d1, extendedExpInc_d2 : std_logic_vector(9 downto 0) := (others => '0');
signal nZerosNew, nZerosNew_d1 : std_logic_vector(4 downto 0) := (others => '0');
signal shiftedFrac, shiftedFrac_d1 : std_logic_vector(27 downto 0) := (others => '0');
signal updatedExp : std_logic_vector(9 downto 0) := (others => '0');
signal eqdiffsign : std_logic := '0';
signal expFrac : std_logic_vector(33 downto 0) := (others => '0');
signal stk : std_logic := '0';
signal rnd : std_logic := '0';
signal grd : std_logic := '0';
signal lsb : std_logic := '0';
signal addToRoundBit, addToRoundBit_d1 : std_logic := '0';
signal RoundedExpFrac : std_logic_vector(33 downto 0) := (others => '0');
signal upExc : std_logic_vector(1 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
signal exExpExc : std_logic_vector(3 downto 0) := (others => '0');
signal excRt2 : std_logic_vector(1 downto 0) := (others => '0');
signal excR : std_logic_vector(1 downto 0) := (others => '0');
signal signR2 : std_logic := '0';
signal computedR : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            newX_d1 <=  newX;
            expX_d1 <=  expX;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            excRt_d1 <=  excRt;
            excRt_d2 <=  excRt_d1;
            excRt_d3 <=  excRt_d2;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            shiftedFracY_d1 <=  shiftedFracY;
            extendedExpInc_d1 <=  extendedExpInc;
            extendedExpInc_d2 <=  extendedExpInc_d1;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            addToRoundBit_d1 <=  addToRoundBit;
         end if;
      end process;
-- Exponent difference and swap  --
   excExpFracX <= X(33 downto 32) & X(30 downto 0);
   excExpFracY <= Y(33 downto 32) & Y(30 downto 0);
   eXmeY <= ("0" & X(30 downto 23)) - ("0" & Y(30 downto 23));
   eYmeX <= ("0" & Y(30 downto 23)) - ("0" & X(30 downto 23));
   swap <= '0' when excExpFracX >= excExpFracY else '1';
   newX <= X when swap = '0' else Y;
   newY <= Y when swap = '0' else X;
   expX<= newX(30 downto 23);
   excX<= newX(33 downto 32);
   excY<= newY(33 downto 32);
   signX<= newX(31);
   signY<= newY(31);
   EffSub <= signX xor signY;
   sXsYExnXY <= signX & signY & excX & excY;
   sdExnXY <= excX & excY;
   fracY <= "000000000000000000000000" when excY="00" else ('1' & newY(22 downto 0));
   with sXsYExnXY select 
   excRt <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR<= '0' when (sXsYExnXY="100000" or sXsYExnXY="010000") else signX;
   ---------------- cycle 0----------------
   expDiff <= eXmeY when swap = '0' else eYmeX;
   shiftedOut <= '1' when (expDiff >= 25) else '0';
   shiftVal <= expDiff(4 downto 0) when shiftedOut='0' else CONV_STD_LOGIC_VECTOR(26,5) ;
   RightShifterComponent: FPAdd_8_23_uid6324686_RightShifter  -- pipelineDepth=0 maxInDelay=2.25704e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal,
                 X => fracY);
   ----------------Synchro barrier, entering cycle 1----------------
   sticky <= '0' when (shiftedFracY_d1(23 downto 0)=CONV_STD_LOGIC_VECTOR(0,23)) else '1';
   ---------------- cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   fracYfar <= "0" & shiftedFracY_d1(49 downto 24);
   EffSubVector <= (26 downto 0 => EffSub_d1);
   fracYfarXorOp <= fracYfar xor EffSubVector;
   fracXfar <= "01" & (newX_d1(22 downto 0)) & "00";
   cInAddFar <= EffSub_d1 and not sticky;
   fracAdder: IntAdder_27_f250_uid6324691  -- pipelineDepth=0 maxInDelay=1.02352e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => cInAddFar,
                 R => fracAddResult,
                 X => fracXfar,
                 Y => fracYfarXorOp);
   fracGRS<= fracAddResult & sticky; 
   extendedExpInc<= ("00" & expX_d1) + '1';
   LZC_component: LZCShifter_28_to_28_counting_32_F250_uid6324698  -- pipelineDepth=1 maxInDelay=1.86552e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => nZerosNew,
                 I => fracGRS,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   updatedExp <= extendedExpInc_d2 - ("00000" & nZerosNew_d1);
   eqdiffsign <= '1' when nZerosNew_d1="11111" else '0';
   expFrac<= updatedExp & shiftedFrac_d1(26 downto 3);
   ---------------- cycle 2----------------
   stk<= shiftedFrac(1) or shiftedFrac(0);
   rnd<= shiftedFrac(2);
   grd<= shiftedFrac(3);
   lsb<= shiftedFrac(4);
   addToRoundBit<= '0' when (lsb='0' and grd='1' and rnd='0' and stk='0')  else '1';
   ----------------Synchro barrier, entering cycle 3----------------
   roundingAdder: IntAdder_34_f250_uid6324701  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => addToRoundBit_d1,
                 R => RoundedExpFrac,
                 X => expFrac,
                 Y => "0000000000000000000000000000000000");
   ---------------- cycle 3----------------
   upExc <= RoundedExpFrac(33 downto 32);
   fracR <= RoundedExpFrac(23 downto 1);
   expR <= RoundedExpFrac(31 downto 24);
   exExpExc <= upExc & excRt_d3;
   with (exExpExc) select 
   excRt2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR <= "00" when (eqdiffsign='1' and EffSub_d3='1') else excRt2;
   signR2 <= '0' when (eqdiffsign='1' and EffSub_d3='1') else signR_d3;
   computedR <= excR & signR2 & expR & fracR;
   R <= computedR;
end architecture;

--------------------------------------------------------------------------------
--         FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          Y : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
   component FPAdd_8_23_uid6324686 is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

signal X_out : std_logic_vector(33 downto 0) := (others => '0');
signal Y_out : std_logic_vector(33 downto 0) := (others => '0');
signal R_temp : std_logic_vector(8+23+2 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
X_out <= X;
Y_out <= Y;
   FPAddSubOp_instance: FPAdd_8_23_uid6324686  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R_temp,
                 X => X_out,
                 Y => Y_out);
   ----------------Synchro barrier, entering cycle 3----------------
R <= R_temp;
end architecture;

--------------------------------------------------------------------------------
--             Mux_sign_1_wordsize_34_numberOfInputs_59_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Mux_sign_1_wordsize_34_numberOfInputs_59_component is
   port ( clk, rst : in std_logic;
          iS_0 : in std_logic_vector(33 downto 0);
          iS_1 : in std_logic_vector(33 downto 0);
          iS_2 : in std_logic_vector(33 downto 0);
          iS_3 : in std_logic_vector(33 downto 0);
          iS_4 : in std_logic_vector(33 downto 0);
          iS_5 : in std_logic_vector(33 downto 0);
          iS_6 : in std_logic_vector(33 downto 0);
          iS_7 : in std_logic_vector(33 downto 0);
          iS_8 : in std_logic_vector(33 downto 0);
          iS_9 : in std_logic_vector(33 downto 0);
          iS_10 : in std_logic_vector(33 downto 0);
          iS_11 : in std_logic_vector(33 downto 0);
          iS_12 : in std_logic_vector(33 downto 0);
          iS_13 : in std_logic_vector(33 downto 0);
          iS_14 : in std_logic_vector(33 downto 0);
          iS_15 : in std_logic_vector(33 downto 0);
          iS_16 : in std_logic_vector(33 downto 0);
          iS_17 : in std_logic_vector(33 downto 0);
          iS_18 : in std_logic_vector(33 downto 0);
          iS_19 : in std_logic_vector(33 downto 0);
          iS_20 : in std_logic_vector(33 downto 0);
          iS_21 : in std_logic_vector(33 downto 0);
          iS_22 : in std_logic_vector(33 downto 0);
          iS_23 : in std_logic_vector(33 downto 0);
          iS_24 : in std_logic_vector(33 downto 0);
          iS_25 : in std_logic_vector(33 downto 0);
          iS_26 : in std_logic_vector(33 downto 0);
          iS_27 : in std_logic_vector(33 downto 0);
          iS_28 : in std_logic_vector(33 downto 0);
          iS_29 : in std_logic_vector(33 downto 0);
          iS_30 : in std_logic_vector(33 downto 0);
          iS_31 : in std_logic_vector(33 downto 0);
          iS_32 : in std_logic_vector(33 downto 0);
          iS_33 : in std_logic_vector(33 downto 0);
          iS_34 : in std_logic_vector(33 downto 0);
          iS_35 : in std_logic_vector(33 downto 0);
          iS_36 : in std_logic_vector(33 downto 0);
          iS_37 : in std_logic_vector(33 downto 0);
          iS_38 : in std_logic_vector(33 downto 0);
          iS_39 : in std_logic_vector(33 downto 0);
          iS_40 : in std_logic_vector(33 downto 0);
          iS_41 : in std_logic_vector(33 downto 0);
          iS_42 : in std_logic_vector(33 downto 0);
          iS_43 : in std_logic_vector(33 downto 0);
          iS_44 : in std_logic_vector(33 downto 0);
          iS_45 : in std_logic_vector(33 downto 0);
          iS_46 : in std_logic_vector(33 downto 0);
          iS_47 : in std_logic_vector(33 downto 0);
          iS_48 : in std_logic_vector(33 downto 0);
          iS_49 : in std_logic_vector(33 downto 0);
          iS_50 : in std_logic_vector(33 downto 0);
          iS_51 : in std_logic_vector(33 downto 0);
          iS_52 : in std_logic_vector(33 downto 0);
          iS_53 : in std_logic_vector(33 downto 0);
          iS_54 : in std_logic_vector(33 downto 0);
          iS_55 : in std_logic_vector(33 downto 0);
          iS_56 : in std_logic_vector(33 downto 0);
          iS_57 : in std_logic_vector(33 downto 0);
          iS_58 : in std_logic_vector(33 downto 0);
          iSel : in std_logic_vector(5 downto 0);
          oMux : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Mux_sign_1_wordsize_34_numberOfInputs_59_component is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   with iSel select
      oMux <= 
         iS_0 when "000000",
         iS_1 when "000001",
         iS_2 when "000010",
         iS_3 when "000011",
         iS_4 when "000100",
         iS_5 when "000101",
         iS_6 when "000110",
         iS_7 when "000111",
         iS_8 when "001000",
         iS_9 when "001001",
         iS_10 when "001010",
         iS_11 when "001011",
         iS_12 when "001100",
         iS_13 when "001101",
         iS_14 when "001110",
         iS_15 when "001111",
         iS_16 when "010000",
         iS_17 when "010001",
         iS_18 when "010010",
         iS_19 when "010011",
         iS_20 when "010100",
         iS_21 when "010101",
         iS_22 when "010110",
         iS_23 when "010111",
         iS_24 when "011000",
         iS_25 when "011001",
         iS_26 when "011010",
         iS_27 when "011011",
         iS_28 when "011100",
         iS_29 when "011101",
         iS_30 when "011110",
         iS_31 when "011111",
         iS_32 when "100000",
         iS_33 when "100001",
         iS_34 when "100010",
         iS_35 when "100011",
         iS_36 when "100100",
         iS_37 when "100101",
         iS_38 when "100110",
         iS_39 when "100111",
         iS_40 when "101000",
         iS_41 when "101001",
         iS_42 when "101010",
         iS_43 when "101011",
         iS_44 when "101100",
         iS_45 when "101101",
         iS_46 when "101110",
         iS_47 when "101111",
         iS_48 when "110000",
         iS_49 when "110001",
         iS_50 when "110010",
         iS_51 when "110011",
         iS_52 when "110100",
         iS_53 when "110101",
         iS_54 when "110110",
         iS_55 when "110111",
         iS_56 when "111000",
         iS_57 when "111001",
         iS_58 when "111010",
(others=>'X') when others;
end architecture;

--------------------------------------------------------------------------------
--                         OutputIEEE_8_23_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. Ferrandi  (2009-2012)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity OutputIEEE_8_23_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(8+23+2 downto 0);
          R : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_component is
signal expX : std_logic_vector(7 downto 0) := (others => '0');
signal fracX : std_logic_vector(22 downto 0) := (others => '0');
signal exnX : std_logic_vector(1 downto 0) := (others => '0');
signal sX : std_logic := '0';
signal expZero : std_logic := '0';
signal sfracX : std_logic_vector(22 downto 0) := (others => '0');
signal fracR : std_logic_vector(22 downto 0) := (others => '0');
signal expR : std_logic_vector(7 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   exnX  <= X(33 downto 32);
   sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
   fracR <= sfracX;
   expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
   R <= sX & expR & fracR; 
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 15 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      Y <= s14;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 16 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      Y <= s15;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 29 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      Y <= s28;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      Y <= s5;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      Y <= s3;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "100100" when "000000",
      "101100" when "000001",
      "100110" when "000010",
      "000111" when "000011",
      "011101" when "000100",
      "010101" when "000101",
      "011010" when "000110",
      "000000" when "000111",
      "001000" when "001000",
      "010010" when "001001",
      "000000" when "001010",
      "011000" when "001011",
      "001100" when "001100",
      "000101" when "001101",
      "011110" when "001110",
      "000000" when "001111",
      "101101" when "010000",
      "100101" when "010001",
      "010110" when "010010",
      "001101" when "010011",
      "101111" when "010100",
      "011011" when "010101",
      "000001" when "010110",
      "001001" when "010111",
      "011111" when "011000",
      "101010" when "011001",
      "011001" when "011010",
      "110010" when "011011",
      "000110" when "011100",
      "100010" when "011101",
      "101110" when "011110",
      "000000" when "011111",
      "110011" when "100000",
      "010111" when "100001",
      "001110" when "100010",
      "110000" when "100011",
      "011100" when "100100",
      "110100" when "100101",
      "010000" when "100110",
      "100000" when "100111",
      "101000" when "101000",
      "001010" when "101001",
      "110101" when "101010",
      "010011" when "101011",
      "100011" when "101100",
      "101011" when "101101",
      "000000" when "101110",
      "110110" when "101111",
      "100111" when "110000",
      "001111" when "110001",
      "110001" when "110010",
      "000010" when "110011",
      "000011" when "110100",
      "010001" when "110101",
      "100001" when "110110",
      "101001" when "110111",
      "001011" when "111000",
      "000100" when "111001",
      "010100" when "111010",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "101100" when "000000",
      "011011" when "000001",
      "000001" when "000010",
      "110000" when "000011",
      "011110" when "000100",
      "001010" when "000101",
      "001101" when "000110",
      "110010" when "000111",
      "001000" when "001000",
      "011001" when "001001",
      "000000" when "001010",
      "110101" when "001011",
      "010010" when "001100",
      "101110" when "001101",
      "011111" when "001110",
      "000000" when "001111",
      "011100" when "010000",
      "000000" when "010001",
      "001011" when "010010",
      "010100" when "010011",
      "000010" when "010100",
      "001110" when "010101",
      "110011" when "010110",
      "001001" when "010111",
      "100111" when "011000",
      "100101" when "011001",
      "110110" when "011010",
      "000101" when "011011",
      "101111" when "011100",
      "101010" when "011101",
      "011101" when "011110",
      "000000" when "011111",
      "000110" when "100000",
      "001100" when "100001",
      "010101" when "100010",
      "000011" when "100011",
      "001111" when "100100",
      "110001" when "100101",
      "010111" when "100110",
      "101000" when "100111",
      "100011" when "101000",
      "010000" when "101001",
      "000111" when "101010",
      "100000" when "101011",
      "101011" when "101100",
      "011010" when "101101",
      "000000" when "101110",
      "010011" when "101111",
      "100010" when "110000",
      "010110" when "110001",
      "000100" when "110010",
      "110100" when "110011",
      "100110" when "110100",
      "011000" when "110101",
      "101001" when "110110",
      "100100" when "110111",
      "010001" when "111000",
      "101101" when "111001",
      "100001" when "111010",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000000" when "000000",
      "000000" when "000001",
      "000000" when "000010",
      "101000" when "000011",
      "011101" when "000100",
      "011111" when "000101",
      "010010" when "000110",
      "000001" when "000111",
      "000100" when "001000",
      "011011" when "001001",
      "000000" when "001010",
      "011110" when "001011",
      "100001" when "001100",
      "100110" when "001101",
      "001010" when "001110",
      "000000" when "001111",
      "000000" when "010000",
      "100011" when "010001",
      "000110" when "010010",
      "011000" when "010011",
      "001100" when "010100",
      "010011" when "010101",
      "000010" when "010110",
      "000101" when "010111",
      "000000" when "011000",
      "000000" when "011001",
      "001001" when "011010",
      "100111" when "011011",
      "001011" when "011100",
      "010101" when "011101",
      "000000" when "011110",
      "000000" when "011111",
      "011100" when "100000",
      "000111" when "100001",
      "011001" when "100010",
      "001101" when "100011",
      "010100" when "100100",
      "000000" when "100101",
      "001000" when "100110",
      "000000" when "100111",
      "000000" when "101000",
      "001111" when "101001",
      "100000" when "101010",
      "000000" when "101011",
      "010110" when "101100",
      "000000" when "101101",
      "000000" when "101110",
      "100010" when "101111",
      "001110" when "110000",
      "011010" when "110001",
      "010001" when "110010",
      "000011" when "110011",
      "100100" when "110100",
      "000000" when "110101",
      "000000" when "110110",
      "010000" when "110111",
      "000000" when "111000",
      "100101" when "111001",
      "010111" when "111010",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--          GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic;
          o5 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(5 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000000" when "000000",
      "000000" when "000001",
      "000000" when "000010",
      "010000" when "000011",
      "011000" when "000100",
      "000010" when "000101",
      "010001" when "000110",
      "100100" when "000111",
      "011101" when "001000",
      "011111" when "001001",
      "000000" when "001010",
      "011001" when "001011",
      "000100" when "001100",
      "001000" when "001101",
      "010110" when "001110",
      "000000" when "001111",
      "000000" when "010000",
      "000110" when "010001",
      "100000" when "010010",
      "011010" when "010011",
      "001011" when "010100",
      "010010" when "010101",
      "100101" when "010110",
      "011110" when "010111",
      "000000" when "011000",
      "000000" when "011001",
      "001111" when "011010",
      "001001" when "011011",
      "010111" when "011100",
      "010100" when "011101",
      "000000" when "011110",
      "000000" when "011111",
      "000001" when "100000",
      "100001" when "100001",
      "011011" when "100010",
      "001100" when "100011",
      "010011" when "100100",
      "100011" when "100101",
      "001010" when "100110",
      "000000" when "100111",
      "000000" when "101000",
      "100111" when "101001",
      "000011" when "101010",
      "000000" when "101011",
      "010101" when "101100",
      "000000" when "101101",
      "000000" when "101110",
      "000101" when "101111",
      "001101" when "110000",
      "011100" when "110001",
      "001110" when "110010",
      "100110" when "110011",
      "100010" when "110100",
      "000000" when "110101",
      "000000" when "110110",
      "101000" when "110111",
      "000000" when "111000",
      "000111" when "111001",
      "000000" when "111010",
      "000000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
   o5 <= t_out(5);
end architecture;

--------------------------------------------------------------------------------
-- GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
   component GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic;
             o5 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
signal Output5_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp,
                 o5 => Output5_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;
Output(5) <= Output5_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "00000" when "000000",
      "00000" when "000001",
      "00000" when "000010",
      "01110" when "000011",
      "00011" when "000100",
      "00000" when "000101",
      "00000" when "000110",
      "00000" when "000111",
      "01111" when "001000",
      "00000" when "001001",
      "00000" when "001010",
      "00000" when "001011",
      "00000" when "001100",
      "00000" when "001101",
      "01010" when "001110",
      "00000" when "001111",
      "00000" when "010000",
      "00000" when "010001",
      "10001" when "010010",
      "00110" when "010011",
      "00000" when "010100",
      "00000" when "010101",
      "10000" when "010110",
      "00100" when "010111",
      "00000" when "011000",
      "00000" when "011001",
      "00000" when "011010",
      "00000" when "011011",
      "00000" when "011100",
      "00000" when "011101",
      "00000" when "011110",
      "00000" when "011111",
      "10010" when "100000",
      "01100" when "100001",
      "00111" when "100010",
      "00000" when "100011",
      "00000" when "100100",
      "00000" when "100101",
      "00000" when "100110",
      "00000" when "100111",
      "00000" when "101000",
      "00000" when "101001",
      "00001" when "101010",
      "00000" when "101011",
      "00000" when "101100",
      "00000" when "101101",
      "00000" when "101110",
      "01011" when "101111",
      "01000" when "110000",
      "00101" when "110001",
      "01001" when "110010",
      "00000" when "110011",
      "00010" when "110100",
      "00000" when "110101",
      "00000" when "110110",
      "00000" when "110111",
      "00000" when "111000",
      "01101" when "111001",
      "00000" when "111010",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic;
          o3 : out std_logic;
          o4 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(4 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "00000" when "000000",
      "00000" when "000001",
      "00000" when "000010",
      "00010" when "000011",
      "00111" when "000100",
      "00000" when "000101",
      "00000" when "000110",
      "00000" when "000111",
      "10000" when "001000",
      "00000" when "001001",
      "00000" when "001010",
      "00000" when "001011",
      "00000" when "001100",
      "00000" when "001101",
      "01110" when "001110",
      "00000" when "001111",
      "00000" when "010000",
      "00000" when "010001",
      "00101" when "010010",
      "01001" when "010011",
      "00000" when "010100",
      "00000" when "010101",
      "10001" when "010110",
      "01000" when "010111",
      "00000" when "011000",
      "00000" when "011001",
      "00000" when "011010",
      "00000" when "011011",
      "00000" when "011100",
      "00000" when "011101",
      "00000" when "011110",
      "00000" when "011111",
      "00110" when "100000",
      "01101" when "100001",
      "01010" when "100010",
      "00000" when "100011",
      "00000" when "100100",
      "10010" when "100101",
      "00000" when "100110",
      "00000" when "100111",
      "00000" when "101000",
      "00000" when "101001",
      "01111" when "101010",
      "00000" when "101011",
      "00000" when "101100",
      "00000" when "101101",
      "00000" when "101110",
      "00000" when "101111",
      "01011" when "110000",
      "00100" when "110001",
      "01100" when "110010",
      "00000" when "110011",
      "00011" when "110100",
      "00000" when "110101",
      "00000" when "110110",
      "00000" when "110111",
      "00000" when "111000",
      "00001" when "111001",
      "00000" when "111010",
      "00000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
   o3 <= t_out(3);
   o4 <= t_out(4);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(4 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5_wrapper_component is
   component GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic;
             o3 : out std_logic;
             o4 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
signal Output3_temp : std_logic := '0';
signal Output4_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp,
                 o3 => Output3_temp,
                 o4 => Output4_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;
Output(3) <= Output3_temp;
Output(4) <= Output4_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product10_3_impl_0_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product10_3_impl_0_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product10_3_impl_0_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "010" when "000011",
      "011" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "100" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "000" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "001" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product10_3_impl_0_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product10_3_impl_0_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product10_3_impl_0_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Product10_3_impl_0_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product10_3_impl_0_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--         GenericLut_LUTData_MUX_Product10_3_impl_1_LUT_wIn_6_wOut_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
-- >> University of Kassel, Germany
-- >> Digital Technology Group
-- >> Author(s):
-- >> Marco Kleinlein <kleinlein@uni-kassel.de>
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product10_3_impl_1_LUT_wIn_6_wOut_3 is
   port ( i0 : in std_logic;
          i1 : in std_logic;
          i2 : in std_logic;
          i3 : in std_logic;
          i4 : in std_logic;
          i5 : in std_logic;
          o0 : out std_logic;
          o1 : out std_logic;
          o2 : out std_logic   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product10_3_impl_1_LUT_wIn_6_wOut_3 is
signal t_in : std_logic_vector(5 downto 0) := (others => '0');
signal t_out : std_logic_vector(2 downto 0) := (others => '0');
begin
   t_in(0) <= i0;
   t_in(1) <= i1;
   t_in(2) <= i2;
   t_in(3) <= i3;
   t_in(4) <= i4;
   t_in(5) <= i5;
   with t_in select t_out <= 
      "000" when "000000",
      "000" when "000001",
      "000" when "000010",
      "000" when "000011",
      "010" when "000100",
      "000" when "000101",
      "000" when "000110",
      "000" when "000111",
      "000" when "001000",
      "000" when "001001",
      "000" when "001010",
      "000" when "001011",
      "000" when "001100",
      "000" when "001101",
      "000" when "001110",
      "000" when "001111",
      "000" when "010000",
      "000" when "010001",
      "000" when "010010",
      "001" when "010011",
      "000" when "010100",
      "000" when "010101",
      "000" when "010110",
      "000" when "010111",
      "000" when "011000",
      "000" when "011001",
      "000" when "011010",
      "000" when "011011",
      "000" when "011100",
      "000" when "011101",
      "000" when "011110",
      "000" when "011111",
      "000" when "100000",
      "000" when "100001",
      "000" when "100010",
      "000" when "100011",
      "000" when "100100",
      "011" when "100101",
      "000" when "100110",
      "000" when "100111",
      "000" when "101000",
      "000" when "101001",
      "000" when "101010",
      "000" when "101011",
      "000" when "101100",
      "000" when "101101",
      "000" when "101110",
      "100" when "101111",
      "000" when "110000",
      "000" when "110001",
      "000" when "110010",
      "000" when "110011",
      "000" when "110100",
      "000" when "110101",
      "000" when "110110",
      "000" when "110111",
      "000" when "111000",
      "000" when "111001",
      "000" when "111010",
      "000" when others;

   o0 <= t_out(0);
   o1 <= t_out(1);
   o2 <= t_out(2);
end architecture;

--------------------------------------------------------------------------------
--GenericLut_LUTData_MUX_Product10_3_impl_1_LUT_wIn_6_wOut_3_wrapper_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity GenericLut_LUTData_MUX_Product10_3_impl_1_LUT_wIn_6_wOut_3_wrapper_component is
   port ( clk, rst : in std_logic;
          Input : in std_logic_vector(5 downto 0);
          Output : out std_logic_vector(2 downto 0)   );
end entity;

architecture arch of GenericLut_LUTData_MUX_Product10_3_impl_1_LUT_wIn_6_wOut_3_wrapper_component is
   component GenericLut_LUTData_MUX_Product10_3_impl_1_LUT_wIn_6_wOut_3 is
      port ( i0 : in std_logic;
             i1 : in std_logic;
             i2 : in std_logic;
             i3 : in std_logic;
             i4 : in std_logic;
             i5 : in std_logic;
             o0 : out std_logic;
             o1 : out std_logic;
             o2 : out std_logic   );
   end component;

signal Input0_out : std_logic := '0';
signal Input1_out : std_logic := '0';
signal Input2_out : std_logic := '0';
signal Input3_out : std_logic := '0';
signal Input4_out : std_logic := '0';
signal Input5_out : std_logic := '0';
signal Output0_temp : std_logic := '0';
signal Output1_temp : std_logic := '0';
signal Output2_temp : std_logic := '0';
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
Input0_out <= Input(0);
Input1_out <= Input(1);
Input2_out <= Input(2);
Input3_out <= Input(3);
Input4_out <= Input(4);
Input5_out <= Input(5);
   instLUT: GenericLut_LUTData_MUX_Product10_3_impl_1_LUT_wIn_6_wOut_3
      port map ( i0 => Input0_out,
                 i1 => Input1_out,
                 i2 => Input2_out,
                 i3 => Input3_out,
                 i4 => Input4_out,
                 i5 => Input5_out,
                 o0 => Output0_temp,
                 o1 => Output1_temp,
                 o2 => Output2_temp);
   ----------------Synchro barrier, entering cycle 0----------------
Output(0) <= Output0_temp;
Output(1) <= Output1_temp;
Output(2) <= Output2_temp;

end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 14 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      Y <= s13;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 20 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      Y <= s19;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 24 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      Y <= s23;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 25 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      Y <= s24;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      Y <= s9;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      Y <= s20;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 28 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      Y <= s27;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      Y <= s2;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 38 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      Y <= s37;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      Y <= s4;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      Y <= s8;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 19 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      Y <= s18;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 35 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      Y <= s34;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 34 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      Y <= s33;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      Y <= s10;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      Y <= s12;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 27 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      Y <= s26;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 26 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      Y <= s25;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 30 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      Y <= s29;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      Y <= s1;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 36 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      Y <= s35;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 37 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      Y <= s36;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      Y <= s7;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      Y <= s6;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 18 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      Y <= s17;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      Y <= s11;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 17 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      Y <= s16;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 23 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      Y <= s22;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 39 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      Y <= s38;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 52 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      Y <= s51;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 57 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      Y <= s56;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 62 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      Y <= s61;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 67 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      Y <= s66;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 41 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      Y <= s40;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_78_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 78 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_78_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_78_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      Y <= s77;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_97_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 97 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_97_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_97_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      Y <= s96;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_102_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 102 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_102_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_102_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      Y <= s101;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 64 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      Y <= s63;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_77_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 77 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_77_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_77_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      Y <= s76;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 65 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      Y <= s64;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_122_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 122 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_122_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_122_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      Y <= s121;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_124_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 124 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_124_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_124_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      Y <= s123;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_132_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 132 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_132_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_132_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      Y <= s131;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_137_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 137 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_137_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_137_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      Y <= s136;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_142_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 142 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_142_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_142_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      Y <= s141;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_147_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 147 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_147_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_147_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
signal s107 : std_logic_vector(33 downto 0) := (others => '0');
signal s108 : std_logic_vector(33 downto 0) := (others => '0');
signal s109 : std_logic_vector(33 downto 0) := (others => '0');
signal s110 : std_logic_vector(33 downto 0) := (others => '0');
signal s111 : std_logic_vector(33 downto 0) := (others => '0');
signal s112 : std_logic_vector(33 downto 0) := (others => '0');
signal s113 : std_logic_vector(33 downto 0) := (others => '0');
signal s114 : std_logic_vector(33 downto 0) := (others => '0');
signal s115 : std_logic_vector(33 downto 0) := (others => '0');
signal s116 : std_logic_vector(33 downto 0) := (others => '0');
signal s117 : std_logic_vector(33 downto 0) := (others => '0');
signal s118 : std_logic_vector(33 downto 0) := (others => '0');
signal s119 : std_logic_vector(33 downto 0) := (others => '0');
signal s120 : std_logic_vector(33 downto 0) := (others => '0');
signal s121 : std_logic_vector(33 downto 0) := (others => '0');
signal s122 : std_logic_vector(33 downto 0) := (others => '0');
signal s123 : std_logic_vector(33 downto 0) := (others => '0');
signal s124 : std_logic_vector(33 downto 0) := (others => '0');
signal s125 : std_logic_vector(33 downto 0) := (others => '0');
signal s126 : std_logic_vector(33 downto 0) := (others => '0');
signal s127 : std_logic_vector(33 downto 0) := (others => '0');
signal s128 : std_logic_vector(33 downto 0) := (others => '0');
signal s129 : std_logic_vector(33 downto 0) := (others => '0');
signal s130 : std_logic_vector(33 downto 0) := (others => '0');
signal s131 : std_logic_vector(33 downto 0) := (others => '0');
signal s132 : std_logic_vector(33 downto 0) := (others => '0');
signal s133 : std_logic_vector(33 downto 0) := (others => '0');
signal s134 : std_logic_vector(33 downto 0) := (others => '0');
signal s135 : std_logic_vector(33 downto 0) := (others => '0');
signal s136 : std_logic_vector(33 downto 0) := (others => '0');
signal s137 : std_logic_vector(33 downto 0) := (others => '0');
signal s138 : std_logic_vector(33 downto 0) := (others => '0');
signal s139 : std_logic_vector(33 downto 0) := (others => '0');
signal s140 : std_logic_vector(33 downto 0) := (others => '0');
signal s141 : std_logic_vector(33 downto 0) := (others => '0');
signal s142 : std_logic_vector(33 downto 0) := (others => '0');
signal s143 : std_logic_vector(33 downto 0) := (others => '0');
signal s144 : std_logic_vector(33 downto 0) := (others => '0');
signal s145 : std_logic_vector(33 downto 0) := (others => '0');
signal s146 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
      s107 <= "0000000000000000000000000000000000";
      s108 <= "0000000000000000000000000000000000";
      s109 <= "0000000000000000000000000000000000";
      s110 <= "0000000000000000000000000000000000";
      s111 <= "0000000000000000000000000000000000";
      s112 <= "0000000000000000000000000000000000";
      s113 <= "0000000000000000000000000000000000";
      s114 <= "0000000000000000000000000000000000";
      s115 <= "0000000000000000000000000000000000";
      s116 <= "0000000000000000000000000000000000";
      s117 <= "0000000000000000000000000000000000";
      s118 <= "0000000000000000000000000000000000";
      s119 <= "0000000000000000000000000000000000";
      s120 <= "0000000000000000000000000000000000";
      s121 <= "0000000000000000000000000000000000";
      s122 <= "0000000000000000000000000000000000";
      s123 <= "0000000000000000000000000000000000";
      s124 <= "0000000000000000000000000000000000";
      s125 <= "0000000000000000000000000000000000";
      s126 <= "0000000000000000000000000000000000";
      s127 <= "0000000000000000000000000000000000";
      s128 <= "0000000000000000000000000000000000";
      s129 <= "0000000000000000000000000000000000";
      s130 <= "0000000000000000000000000000000000";
      s131 <= "0000000000000000000000000000000000";
      s132 <= "0000000000000000000000000000000000";
      s133 <= "0000000000000000000000000000000000";
      s134 <= "0000000000000000000000000000000000";
      s135 <= "0000000000000000000000000000000000";
      s136 <= "0000000000000000000000000000000000";
      s137 <= "0000000000000000000000000000000000";
      s138 <= "0000000000000000000000000000000000";
      s139 <= "0000000000000000000000000000000000";
      s140 <= "0000000000000000000000000000000000";
      s141 <= "0000000000000000000000000000000000";
      s142 <= "0000000000000000000000000000000000";
      s143 <= "0000000000000000000000000000000000";
      s144 <= "0000000000000000000000000000000000";
      s145 <= "0000000000000000000000000000000000";
      s146 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      s107 <= s106;
      s108 <= s107;
      s109 <= s108;
      s110 <= s109;
      s111 <= s110;
      s112 <= s111;
      s113 <= s112;
      s114 <= s113;
      s115 <= s114;
      s116 <= s115;
      s117 <= s116;
      s118 <= s117;
      s119 <= s118;
      s120 <= s119;
      s121 <= s120;
      s122 <= s121;
      s123 <= s122;
      s124 <= s123;
      s125 <= s124;
      s126 <= s125;
      s127 <= s126;
      s128 <= s127;
      s129 <= s128;
      s130 <= s129;
      s131 <= s130;
      s132 <= s131;
      s133 <= s132;
      s134 <= s133;
      s135 <= s134;
      s136 <= s135;
      s137 <= s136;
      s138 <= s137;
      s139 <= s138;
      s140 <= s139;
      s141 <= s140;
      s142 <= s141;
      s143 <= s142;
      s144 <= s143;
      s145 <= s144;
      s146 <= s145;
      Y <= s146;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 107 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
signal s104 : std_logic_vector(33 downto 0) := (others => '0');
signal s105 : std_logic_vector(33 downto 0) := (others => '0');
signal s106 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
      s104 <= "0000000000000000000000000000000000";
      s105 <= "0000000000000000000000000000000000";
      s106 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      s104 <= s103;
      s105 <= s104;
      s106 <= s105;
      Y <= s106;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 99 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      Y <= s98;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_104_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 104 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_104_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_104_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
signal s47 : std_logic_vector(33 downto 0) := (others => '0');
signal s48 : std_logic_vector(33 downto 0) := (others => '0');
signal s49 : std_logic_vector(33 downto 0) := (others => '0');
signal s50 : std_logic_vector(33 downto 0) := (others => '0');
signal s51 : std_logic_vector(33 downto 0) := (others => '0');
signal s52 : std_logic_vector(33 downto 0) := (others => '0');
signal s53 : std_logic_vector(33 downto 0) := (others => '0');
signal s54 : std_logic_vector(33 downto 0) := (others => '0');
signal s55 : std_logic_vector(33 downto 0) := (others => '0');
signal s56 : std_logic_vector(33 downto 0) := (others => '0');
signal s57 : std_logic_vector(33 downto 0) := (others => '0');
signal s58 : std_logic_vector(33 downto 0) := (others => '0');
signal s59 : std_logic_vector(33 downto 0) := (others => '0');
signal s60 : std_logic_vector(33 downto 0) := (others => '0');
signal s61 : std_logic_vector(33 downto 0) := (others => '0');
signal s62 : std_logic_vector(33 downto 0) := (others => '0');
signal s63 : std_logic_vector(33 downto 0) := (others => '0');
signal s64 : std_logic_vector(33 downto 0) := (others => '0');
signal s65 : std_logic_vector(33 downto 0) := (others => '0');
signal s66 : std_logic_vector(33 downto 0) := (others => '0');
signal s67 : std_logic_vector(33 downto 0) := (others => '0');
signal s68 : std_logic_vector(33 downto 0) := (others => '0');
signal s69 : std_logic_vector(33 downto 0) := (others => '0');
signal s70 : std_logic_vector(33 downto 0) := (others => '0');
signal s71 : std_logic_vector(33 downto 0) := (others => '0');
signal s72 : std_logic_vector(33 downto 0) := (others => '0');
signal s73 : std_logic_vector(33 downto 0) := (others => '0');
signal s74 : std_logic_vector(33 downto 0) := (others => '0');
signal s75 : std_logic_vector(33 downto 0) := (others => '0');
signal s76 : std_logic_vector(33 downto 0) := (others => '0');
signal s77 : std_logic_vector(33 downto 0) := (others => '0');
signal s78 : std_logic_vector(33 downto 0) := (others => '0');
signal s79 : std_logic_vector(33 downto 0) := (others => '0');
signal s80 : std_logic_vector(33 downto 0) := (others => '0');
signal s81 : std_logic_vector(33 downto 0) := (others => '0');
signal s82 : std_logic_vector(33 downto 0) := (others => '0');
signal s83 : std_logic_vector(33 downto 0) := (others => '0');
signal s84 : std_logic_vector(33 downto 0) := (others => '0');
signal s85 : std_logic_vector(33 downto 0) := (others => '0');
signal s86 : std_logic_vector(33 downto 0) := (others => '0');
signal s87 : std_logic_vector(33 downto 0) := (others => '0');
signal s88 : std_logic_vector(33 downto 0) := (others => '0');
signal s89 : std_logic_vector(33 downto 0) := (others => '0');
signal s90 : std_logic_vector(33 downto 0) := (others => '0');
signal s91 : std_logic_vector(33 downto 0) := (others => '0');
signal s92 : std_logic_vector(33 downto 0) := (others => '0');
signal s93 : std_logic_vector(33 downto 0) := (others => '0');
signal s94 : std_logic_vector(33 downto 0) := (others => '0');
signal s95 : std_logic_vector(33 downto 0) := (others => '0');
signal s96 : std_logic_vector(33 downto 0) := (others => '0');
signal s97 : std_logic_vector(33 downto 0) := (others => '0');
signal s98 : std_logic_vector(33 downto 0) := (others => '0');
signal s99 : std_logic_vector(33 downto 0) := (others => '0');
signal s100 : std_logic_vector(33 downto 0) := (others => '0');
signal s101 : std_logic_vector(33 downto 0) := (others => '0');
signal s102 : std_logic_vector(33 downto 0) := (others => '0');
signal s103 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
      s47 <= "0000000000000000000000000000000000";
      s48 <= "0000000000000000000000000000000000";
      s49 <= "0000000000000000000000000000000000";
      s50 <= "0000000000000000000000000000000000";
      s51 <= "0000000000000000000000000000000000";
      s52 <= "0000000000000000000000000000000000";
      s53 <= "0000000000000000000000000000000000";
      s54 <= "0000000000000000000000000000000000";
      s55 <= "0000000000000000000000000000000000";
      s56 <= "0000000000000000000000000000000000";
      s57 <= "0000000000000000000000000000000000";
      s58 <= "0000000000000000000000000000000000";
      s59 <= "0000000000000000000000000000000000";
      s60 <= "0000000000000000000000000000000000";
      s61 <= "0000000000000000000000000000000000";
      s62 <= "0000000000000000000000000000000000";
      s63 <= "0000000000000000000000000000000000";
      s64 <= "0000000000000000000000000000000000";
      s65 <= "0000000000000000000000000000000000";
      s66 <= "0000000000000000000000000000000000";
      s67 <= "0000000000000000000000000000000000";
      s68 <= "0000000000000000000000000000000000";
      s69 <= "0000000000000000000000000000000000";
      s70 <= "0000000000000000000000000000000000";
      s71 <= "0000000000000000000000000000000000";
      s72 <= "0000000000000000000000000000000000";
      s73 <= "0000000000000000000000000000000000";
      s74 <= "0000000000000000000000000000000000";
      s75 <= "0000000000000000000000000000000000";
      s76 <= "0000000000000000000000000000000000";
      s77 <= "0000000000000000000000000000000000";
      s78 <= "0000000000000000000000000000000000";
      s79 <= "0000000000000000000000000000000000";
      s80 <= "0000000000000000000000000000000000";
      s81 <= "0000000000000000000000000000000000";
      s82 <= "0000000000000000000000000000000000";
      s83 <= "0000000000000000000000000000000000";
      s84 <= "0000000000000000000000000000000000";
      s85 <= "0000000000000000000000000000000000";
      s86 <= "0000000000000000000000000000000000";
      s87 <= "0000000000000000000000000000000000";
      s88 <= "0000000000000000000000000000000000";
      s89 <= "0000000000000000000000000000000000";
      s90 <= "0000000000000000000000000000000000";
      s91 <= "0000000000000000000000000000000000";
      s92 <= "0000000000000000000000000000000000";
      s93 <= "0000000000000000000000000000000000";
      s94 <= "0000000000000000000000000000000000";
      s95 <= "0000000000000000000000000000000000";
      s96 <= "0000000000000000000000000000000000";
      s97 <= "0000000000000000000000000000000000";
      s98 <= "0000000000000000000000000000000000";
      s99 <= "0000000000000000000000000000000000";
      s100 <= "0000000000000000000000000000000000";
      s101 <= "0000000000000000000000000000000000";
      s102 <= "0000000000000000000000000000000000";
      s103 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      s47 <= s46;
      s48 <= s47;
      s49 <= s48;
      s50 <= s49;
      s51 <= s50;
      s52 <= s51;
      s53 <= s52;
      s54 <= s53;
      s55 <= s54;
      s56 <= s55;
      s57 <= s56;
      s58 <= s57;
      s59 <= s58;
      s60 <= s59;
      s61 <= s60;
      s62 <= s61;
      s63 <= s62;
      s64 <= s63;
      s65 <= s64;
      s66 <= s65;
      s67 <= s66;
      s68 <= s67;
      s69 <= s68;
      s70 <= s69;
      s71 <= s70;
      s72 <= s71;
      s73 <= s72;
      s74 <= s73;
      s75 <= s74;
      s76 <= s75;
      s77 <= s76;
      s78 <= s77;
      s79 <= s78;
      s80 <= s79;
      s81 <= s80;
      s82 <= s81;
      s83 <= s82;
      s84 <= s83;
      s85 <= s84;
      s86 <= s85;
      s87 <= s86;
      s88 <= s87;
      s89 <= s88;
      s90 <= s89;
      s91 <= s90;
      s92 <= s91;
      s93 <= s92;
      s94 <= s93;
      s95 <= s94;
      s96 <= s95;
      s97 <= s96;
      s98 <= s97;
      s99 <= s98;
      s100 <= s99;
      s101 <= s100;
      s102 <= s101;
      s103 <= s102;
      Y <= s103;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 32 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      Y <= s31;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 42 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      Y <= s41;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Nigel Kretschmer
--------------------------------------------------------------------------------
-- Pipeline depth: 47 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
   port ( clk, rst : in std_logic;
          X : in std_logic_vector(33 downto 0);
          Y : out std_logic_vector(33 downto 0)   );
end entity;

architecture arch of Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
signal s0 : std_logic_vector(33 downto 0) := (others => '0');
signal s1 : std_logic_vector(33 downto 0) := (others => '0');
signal s2 : std_logic_vector(33 downto 0) := (others => '0');
signal s3 : std_logic_vector(33 downto 0) := (others => '0');
signal s4 : std_logic_vector(33 downto 0) := (others => '0');
signal s5 : std_logic_vector(33 downto 0) := (others => '0');
signal s6 : std_logic_vector(33 downto 0) := (others => '0');
signal s7 : std_logic_vector(33 downto 0) := (others => '0');
signal s8 : std_logic_vector(33 downto 0) := (others => '0');
signal s9 : std_logic_vector(33 downto 0) := (others => '0');
signal s10 : std_logic_vector(33 downto 0) := (others => '0');
signal s11 : std_logic_vector(33 downto 0) := (others => '0');
signal s12 : std_logic_vector(33 downto 0) := (others => '0');
signal s13 : std_logic_vector(33 downto 0) := (others => '0');
signal s14 : std_logic_vector(33 downto 0) := (others => '0');
signal s15 : std_logic_vector(33 downto 0) := (others => '0');
signal s16 : std_logic_vector(33 downto 0) := (others => '0');
signal s17 : std_logic_vector(33 downto 0) := (others => '0');
signal s18 : std_logic_vector(33 downto 0) := (others => '0');
signal s19 : std_logic_vector(33 downto 0) := (others => '0');
signal s20 : std_logic_vector(33 downto 0) := (others => '0');
signal s21 : std_logic_vector(33 downto 0) := (others => '0');
signal s22 : std_logic_vector(33 downto 0) := (others => '0');
signal s23 : std_logic_vector(33 downto 0) := (others => '0');
signal s24 : std_logic_vector(33 downto 0) := (others => '0');
signal s25 : std_logic_vector(33 downto 0) := (others => '0');
signal s26 : std_logic_vector(33 downto 0) := (others => '0');
signal s27 : std_logic_vector(33 downto 0) := (others => '0');
signal s28 : std_logic_vector(33 downto 0) := (others => '0');
signal s29 : std_logic_vector(33 downto 0) := (others => '0');
signal s30 : std_logic_vector(33 downto 0) := (others => '0');
signal s31 : std_logic_vector(33 downto 0) := (others => '0');
signal s32 : std_logic_vector(33 downto 0) := (others => '0');
signal s33 : std_logic_vector(33 downto 0) := (others => '0');
signal s34 : std_logic_vector(33 downto 0) := (others => '0');
signal s35 : std_logic_vector(33 downto 0) := (others => '0');
signal s36 : std_logic_vector(33 downto 0) := (others => '0');
signal s37 : std_logic_vector(33 downto 0) := (others => '0');
signal s38 : std_logic_vector(33 downto 0) := (others => '0');
signal s39 : std_logic_vector(33 downto 0) := (others => '0');
signal s40 : std_logic_vector(33 downto 0) := (others => '0');
signal s41 : std_logic_vector(33 downto 0) := (others => '0');
signal s42 : std_logic_vector(33 downto 0) := (others => '0');
signal s43 : std_logic_vector(33 downto 0) := (others => '0');
signal s44 : std_logic_vector(33 downto 0) := (others => '0');
signal s45 : std_logic_vector(33 downto 0) := (others => '0');
signal s46 : std_logic_vector(33 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
process(clk, rst, X)
begin
   if rst = '1' then
      Y <= "0000000000000000000000000000000000";
      s1 <= "0000000000000000000000000000000000";
      s2 <= "0000000000000000000000000000000000";
      s3 <= "0000000000000000000000000000000000";
      s4 <= "0000000000000000000000000000000000";
      s5 <= "0000000000000000000000000000000000";
      s6 <= "0000000000000000000000000000000000";
      s7 <= "0000000000000000000000000000000000";
      s8 <= "0000000000000000000000000000000000";
      s9 <= "0000000000000000000000000000000000";
      s10 <= "0000000000000000000000000000000000";
      s11 <= "0000000000000000000000000000000000";
      s12 <= "0000000000000000000000000000000000";
      s13 <= "0000000000000000000000000000000000";
      s14 <= "0000000000000000000000000000000000";
      s15 <= "0000000000000000000000000000000000";
      s16 <= "0000000000000000000000000000000000";
      s17 <= "0000000000000000000000000000000000";
      s18 <= "0000000000000000000000000000000000";
      s19 <= "0000000000000000000000000000000000";
      s20 <= "0000000000000000000000000000000000";
      s21 <= "0000000000000000000000000000000000";
      s22 <= "0000000000000000000000000000000000";
      s23 <= "0000000000000000000000000000000000";
      s24 <= "0000000000000000000000000000000000";
      s25 <= "0000000000000000000000000000000000";
      s26 <= "0000000000000000000000000000000000";
      s27 <= "0000000000000000000000000000000000";
      s28 <= "0000000000000000000000000000000000";
      s29 <= "0000000000000000000000000000000000";
      s30 <= "0000000000000000000000000000000000";
      s31 <= "0000000000000000000000000000000000";
      s32 <= "0000000000000000000000000000000000";
      s33 <= "0000000000000000000000000000000000";
      s34 <= "0000000000000000000000000000000000";
      s35 <= "0000000000000000000000000000000000";
      s36 <= "0000000000000000000000000000000000";
      s37 <= "0000000000000000000000000000000000";
      s38 <= "0000000000000000000000000000000000";
      s39 <= "0000000000000000000000000000000000";
      s40 <= "0000000000000000000000000000000000";
      s41 <= "0000000000000000000000000000000000";
      s42 <= "0000000000000000000000000000000000";
      s43 <= "0000000000000000000000000000000000";
      s44 <= "0000000000000000000000000000000000";
      s45 <= "0000000000000000000000000000000000";
      s46 <= "0000000000000000000000000000000000";
   elsif rising_edge(clk) then
      s1 <= s0;
      s2 <= s1;
      s3 <= s2;
      s4 <= s3;
      s5 <= s4;
      s6 <= s5;
      s7 <= s6;
      s8 <= s7;
      s9 <= s8;
      s10 <= s9;
      s11 <= s10;
      s12 <= s11;
      s13 <= s12;
      s14 <= s13;
      s15 <= s14;
      s16 <= s15;
      s17 <= s16;
      s18 <= s17;
      s19 <= s18;
      s20 <= s19;
      s21 <= s20;
      s22 <= s21;
      s23 <= s22;
      s24 <= s23;
      s25 <= s24;
      s26 <= s25;
      s27 <= s26;
      s28 <= s27;
      s29 <= s28;
      s30 <= s29;
      s31 <= s30;
      s32 <= s31;
      s33 <= s32;
      s34 <= s33;
      s35 <= s34;
      s36 <= s35;
      s37 <= s36;
      s38 <= s37;
      s39 <= s38;
      s40 <= s39;
      s41 <= s40;
      s42 <= s41;
      s43 <= s42;
      s44 <= s43;
      s45 <= s44;
      s46 <= s45;
      Y <= s46;
   end if;
   s0 <= X;
end process;
end architecture;

--------------------------------------------------------------------------------
--                         implementedSystem_toplevel
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity implementedSystem_toplevel is
   port ( clk, rst : in std_logic;
          X_0 : in std_logic_vector(31 downto 0);
          X_1 : in std_logic_vector(31 downto 0);
          X_2 : in std_logic_vector(31 downto 0);
          X_3 : in std_logic_vector(31 downto 0);
          Y_0 : out std_logic_vector(31 downto 0);
          Y_1 : out std_logic_vector(31 downto 0);
          Y_2 : out std_logic_vector(31 downto 0);
          Y_3 : out std_logic_vector(31 downto 0)   );
end entity;

architecture arch of implementedSystem_toplevel is
   component ModuloCounter_59_component is
      port ( clk, rst : in std_logic;
             Counter_out : out std_logic_vector(5 downto 0)   );
   end component;

   component InputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(31 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_31_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_28_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n352_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n432_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n500_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n532_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n129_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_158_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_526_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_964_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n529_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n464_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_29_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n336_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_3136_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_3648_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_4110_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_4478_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_4737_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_4868_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_22_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_1472_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_2008_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_2576_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_8_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n17_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n59_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n116_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n188_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Constant_float_8_23_n268_div_65536_component is
      port ( clk, rst : in std_logic;
             Y : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_55_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iS_47 : in std_logic_vector(33 downto 0);
             iS_48 : in std_logic_vector(33 downto 0);
             iS_49 : in std_logic_vector(33 downto 0);
             iS_50 : in std_logic_vector(33 downto 0);
             iS_51 : in std_logic_vector(33 downto 0);
             iS_52 : in std_logic_vector(33 downto 0);
             iS_53 : in std_logic_vector(33 downto 0);
             iS_54 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_41_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_19_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(4 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_5_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(2 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             Y : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(8+23+2 downto 0)   );
   end component;

   component Mux_sign_1_wordsize_34_numberOfInputs_59_component is
      port ( clk, rst : in std_logic;
             iS_0 : in std_logic_vector(33 downto 0);
             iS_1 : in std_logic_vector(33 downto 0);
             iS_2 : in std_logic_vector(33 downto 0);
             iS_3 : in std_logic_vector(33 downto 0);
             iS_4 : in std_logic_vector(33 downto 0);
             iS_5 : in std_logic_vector(33 downto 0);
             iS_6 : in std_logic_vector(33 downto 0);
             iS_7 : in std_logic_vector(33 downto 0);
             iS_8 : in std_logic_vector(33 downto 0);
             iS_9 : in std_logic_vector(33 downto 0);
             iS_10 : in std_logic_vector(33 downto 0);
             iS_11 : in std_logic_vector(33 downto 0);
             iS_12 : in std_logic_vector(33 downto 0);
             iS_13 : in std_logic_vector(33 downto 0);
             iS_14 : in std_logic_vector(33 downto 0);
             iS_15 : in std_logic_vector(33 downto 0);
             iS_16 : in std_logic_vector(33 downto 0);
             iS_17 : in std_logic_vector(33 downto 0);
             iS_18 : in std_logic_vector(33 downto 0);
             iS_19 : in std_logic_vector(33 downto 0);
             iS_20 : in std_logic_vector(33 downto 0);
             iS_21 : in std_logic_vector(33 downto 0);
             iS_22 : in std_logic_vector(33 downto 0);
             iS_23 : in std_logic_vector(33 downto 0);
             iS_24 : in std_logic_vector(33 downto 0);
             iS_25 : in std_logic_vector(33 downto 0);
             iS_26 : in std_logic_vector(33 downto 0);
             iS_27 : in std_logic_vector(33 downto 0);
             iS_28 : in std_logic_vector(33 downto 0);
             iS_29 : in std_logic_vector(33 downto 0);
             iS_30 : in std_logic_vector(33 downto 0);
             iS_31 : in std_logic_vector(33 downto 0);
             iS_32 : in std_logic_vector(33 downto 0);
             iS_33 : in std_logic_vector(33 downto 0);
             iS_34 : in std_logic_vector(33 downto 0);
             iS_35 : in std_logic_vector(33 downto 0);
             iS_36 : in std_logic_vector(33 downto 0);
             iS_37 : in std_logic_vector(33 downto 0);
             iS_38 : in std_logic_vector(33 downto 0);
             iS_39 : in std_logic_vector(33 downto 0);
             iS_40 : in std_logic_vector(33 downto 0);
             iS_41 : in std_logic_vector(33 downto 0);
             iS_42 : in std_logic_vector(33 downto 0);
             iS_43 : in std_logic_vector(33 downto 0);
             iS_44 : in std_logic_vector(33 downto 0);
             iS_45 : in std_logic_vector(33 downto 0);
             iS_46 : in std_logic_vector(33 downto 0);
             iS_47 : in std_logic_vector(33 downto 0);
             iS_48 : in std_logic_vector(33 downto 0);
             iS_49 : in std_logic_vector(33 downto 0);
             iS_50 : in std_logic_vector(33 downto 0);
             iS_51 : in std_logic_vector(33 downto 0);
             iS_52 : in std_logic_vector(33 downto 0);
             iS_53 : in std_logic_vector(33 downto 0);
             iS_54 : in std_logic_vector(33 downto 0);
             iS_55 : in std_logic_vector(33 downto 0);
             iS_56 : in std_logic_vector(33 downto 0);
             iS_57 : in std_logic_vector(33 downto 0);
             iS_58 : in std_logic_vector(33 downto 0);
             iSel : in std_logic_vector(5 downto 0);
             oMux : out std_logic_vector(33 downto 0)   );
   end component;

   component OutputIEEE_8_23_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(8+23+2 downto 0);
             R : out std_logic_vector(31 downto 0)   );
   end component;

   component Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(5 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(4 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product10_3_impl_0_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component GenericLut_LUTData_MUX_Product10_3_impl_1_LUT_wIn_6_wOut_3_wrapper_component is
      port ( clk, rst : in std_logic;
             Input : in std_logic_vector(5 downto 0);
             Output : out std_logic_vector(2 downto 0)   );
   end component;

   component Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_78_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_97_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_102_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_77_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_122_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_124_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_132_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_137_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_142_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_147_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_104_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

   component Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component is
      port ( clk, rst : in std_logic;
             X : in std_logic_vector(33 downto 0);
             Y : out std_logic_vector(33 downto 0)   );
   end component;

signal ModCount591_out : std_logic_vector(5 downto 0) := (others => '0');
signal X_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal X_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal X_2_out : std_logic_vector(33 downto 0) := (others => '0');
signal X_3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant1_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant10_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant11_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant12_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant13_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant14_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant15_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant16_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant17_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant18_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant19_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant2_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant20_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant21_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant22_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant23_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant24_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant25_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant29_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant3_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant32_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant33_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant34_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant4_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant5_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant6_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant7_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant8_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Constant9_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product1_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product1_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product1_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out : std_logic_vector(33 downto 0) := (others => '0');
signal Product10_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product10_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product10_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Sum10_0_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum10_0_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum10_0_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out : std_logic_vector(33 downto 0) := (others => '0');
signal Sum10_1_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum10_1_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum10_1_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out : std_logic_vector(33 downto 0) := (others => '0');
signal Sum10_2_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum10_2_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum10_2_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out : std_logic_vector(33 downto 0) := (others => '0');
signal Sum10_3_impl_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum10_3_impl_0_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Sum10_3_impl_1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No16_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No17_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No18_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No19_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay871No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay871No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay871No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay872No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay47No7_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No6_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay123No_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay123No1_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay123No2_out : std_logic_vector(33 downto 0) := (others => '0');
signal Delay123No3_out : std_logic_vector(33 downto 0) := (others => '0');
signal MUX_Product_0_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product_0_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product_2_impl_0_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product_2_impl_1_LUT_out : std_logic_vector(5 downto 0) := (others => '0');
signal MUX_Product1_2_impl_0_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal MUX_Product1_2_impl_1_LUT_out : std_logic_vector(4 downto 0) := (others => '0');
signal MUX_Product10_3_impl_0_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal MUX_Product10_3_impl_1_LUT_out : std_logic_vector(2 downto 0) := (others => '0');
signal SharedReg_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out : std_logic_vector(33 downto 0) := (others => '0');
signal X_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal X_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal X_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal X_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Delay1No_out_to_Product_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No1_out_to_Product_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg249_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg285_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg286_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg279_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg283_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg284_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg305_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg326_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg287_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg308_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg329_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg292_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg290_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg289_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg310_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg288_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg291_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg312_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg354_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg282_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg295_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg316_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg337_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg293_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg314_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg335_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg278_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg280_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg281_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg276_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg297_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No2_out_to_Product_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No3_out_to_Product_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg226_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg232_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg235_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg238_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg239_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg242_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg244_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg248_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg250_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg254_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg353_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg300_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg307_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg299_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg320_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg306_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg327_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg342_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg304_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg294_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg315_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg336_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg311_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg332_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg331_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg352_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg309_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg333_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay123No_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay123No1_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay123No2_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg303_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg324_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg358_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg301_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg322_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg302_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg277_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg298_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg340_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg318_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg339_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No4_out_to_Product1_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No5_out_to_Product1_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg227_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg229_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg231_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg233_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg234_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg236_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg240_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg241_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg245_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg246_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg251_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg252_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg253_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg255_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg321_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg328_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg348_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg325_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg346_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg347_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg350_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg313_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg334_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg355_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg357_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg351_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg356_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg341_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg323_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg344_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg319_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No6_out_to_Product10_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No7_out_to_Product10_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg228_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg230_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg237_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg243_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg247_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg349_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg330_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay123No3_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg345_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg343_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No8_out_to_Sum10_0_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No9_out_to_Sum10_0_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg170_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg191_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg114_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg59_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg118_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg80_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg133_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg4_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg25_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg174_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg63_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg178_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg8_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg122_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg19_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg73_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg126_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg197_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg190_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg67_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg12_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg139_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg71_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg182_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg131_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg168_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay871No1_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg144_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg224_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg53_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg29_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg204_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg108_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg259_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg84_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg164_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg89_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg160_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg152_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg105_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg217_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg93_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg38_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg35_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg213_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg143_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg97_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg149_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg46_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg101_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg202_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg42_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg157_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg210_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No10_out_to_Sum10_1_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No11_out_to_Sum10_1_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg27_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg21_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg123_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg68_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg196_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg127_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg13_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg187_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg1_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg56_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg22_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg171_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg115_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg175_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg137_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg189_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg60_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg81_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg5_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg119_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg79_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg9_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg16_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg64_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg179_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg75_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg130_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg183_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg200_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg154_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg206_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg102_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg158_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg32_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg98_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg214_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg40_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg225_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay871No2_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg201_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg54_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg109_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg50_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg85_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg34_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg165_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg257_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg141_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg221_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg146_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg218_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg209_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg161_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg47_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg150_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg94_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg91_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg43_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No12_out_to_Sum10_2_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No13_out_to_Sum10_2_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg65_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg72_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg120_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg10_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg132_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg186_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg193_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg14_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg83_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg129_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg77_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg180_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg124_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg26_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg184_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg69_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg18_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg57_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg112_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg78_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg2_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg172_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg6_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg194_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg20_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg116_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg138_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg61_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg176_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg136_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg48_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg39_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg263_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg219_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg103_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg261_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg207_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg151_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg148_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg99_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg30_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg211_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg36_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg215_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg88_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg155_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg44_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg269_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg96_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg55_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay872No_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg31_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg110_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg166_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg106_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg142_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg267_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg90_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg222_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg268_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg198_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg51_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg163_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg203_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg258_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg262_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No14_out_to_Sum10_3_impl_parent_implementedSystem_port_0_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay1No15_out_to_Sum10_3_impl_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg173_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg195_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg117_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg7_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg192_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg121_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg128_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg177_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg66_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg188_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg17_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg23_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg70_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg140_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg185_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg134_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg11_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg181_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg82_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg15_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg125_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg74_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg113_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg169_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg135_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg58_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg3_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg62_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg24_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg76_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg52_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_1_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg265_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_2_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg273_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_3_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_4_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg28_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_5_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg107_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_6_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg256_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_7_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_8_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_9_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg220_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_10_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg33_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_11_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg266_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_12_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg270_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_13_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_14_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg104_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_15_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg95_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_16_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_17_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay47No7_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_18_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_19_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg49_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_20_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg159_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_21_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_22_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay15No6_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_23_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg37_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_24_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg208_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_25_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg205_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_26_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_27_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_28_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg156_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_29_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg86_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_30_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg41_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_31_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_32_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_33_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg92_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_34_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg216_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_35_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg45_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_36_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_37_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_38_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg145_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_39_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg212_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_40_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg100_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_41_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_42_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_43_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg153_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_44_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg111_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_45_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Delay871No_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_46_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_47_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg260_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_48_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg87_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_49_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg167_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_50_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg223_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_51_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg274_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_52_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_53_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg162_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_54_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg199_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_55_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_56_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_57_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg272_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_58_cast : std_logic_vector(33 downto 0) := (others => '0');
signal SharedReg147_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_59_cast : std_logic_vector(33 downto 0) := (others => '0');
signal Y_0_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Y_1_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Y_2_IEEE : std_logic_vector(31 downto 0) := (others => '0');
signal Y_3_IEEE : std_logic_vector(31 downto 0) := (others => '0');
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   ModCount591_instance: ModuloCounter_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Counter_out => ModCount591_out);
X_0_IEEE <= X_0;
   X_0_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => X_0_out,
                 X => X_0_IEEE);
X_1_IEEE <= X_1;
   X_1_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => X_1_out,
                 X => X_1_IEEE);
X_2_IEEE <= X_2;
   X_2_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => X_2_out,
                 X => X_2_IEEE);
X_3_IEEE <= X_3;
   X_3_instance: InputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => X_3_out,
                 X => X_3_IEEE);
   Constant_0_impl_instance: Constant_float_8_23_31_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant_0_impl_out);
   Constant1_0_impl_instance: Constant_float_8_23_28_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant1_0_impl_out);
   Constant10_0_impl_instance: Constant_float_8_23_n352_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant10_0_impl_out);
   Constant11_0_impl_instance: Constant_float_8_23_n432_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant11_0_impl_out);
   Constant12_0_impl_instance: Constant_float_8_23_n500_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant12_0_impl_out);
   Constant13_0_impl_instance: Constant_float_8_23_n532_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant13_0_impl_out);
   Constant14_0_impl_instance: Constant_float_8_23_n129_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant14_0_impl_out);
   Constant15_0_impl_instance: Constant_float_8_23_158_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant15_0_impl_out);
   Constant16_0_impl_instance: Constant_float_8_23_526_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant16_0_impl_out);
   Constant17_0_impl_instance: Constant_float_8_23_964_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant17_0_impl_out);
   Constant18_0_impl_instance: Constant_float_8_23_n529_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant18_0_impl_out);
   Constant19_0_impl_instance: Constant_float_8_23_n464_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant19_0_impl_out);
   Constant2_0_impl_instance: Constant_float_8_23_29_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant2_0_impl_out);
   Constant20_0_impl_instance: Constant_float_8_23_n336_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant20_0_impl_out);
   Constant21_0_impl_instance: Constant_float_8_23_3136_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant21_0_impl_out);
   Constant22_0_impl_instance: Constant_float_8_23_3648_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant22_0_impl_out);
   Constant23_0_impl_instance: Constant_float_8_23_4110_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant23_0_impl_out);
   Constant24_0_impl_instance: Constant_float_8_23_4478_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant24_0_impl_out);
   Constant25_0_impl_instance: Constant_float_8_23_4737_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant25_0_impl_out);
   Constant29_0_impl_instance: Constant_float_8_23_4868_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant29_0_impl_out);
   Constant3_0_impl_instance: Constant_float_8_23_22_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant3_0_impl_out);
   Constant32_0_impl_instance: Constant_float_8_23_1472_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant32_0_impl_out);
   Constant33_0_impl_instance: Constant_float_8_23_2008_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant33_0_impl_out);
   Constant34_0_impl_instance: Constant_float_8_23_2576_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant34_0_impl_out);
   Constant4_0_impl_instance: Constant_float_8_23_8_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant4_0_impl_out);
   Constant5_0_impl_instance: Constant_float_8_23_n17_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant5_0_impl_out);
   Constant6_0_impl_instance: Constant_float_8_23_n59_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant6_0_impl_out);
   Constant7_0_impl_instance: Constant_float_8_23_n116_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant7_0_impl_out);
   Constant8_0_impl_instance: Constant_float_8_23_n188_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant8_0_impl_out);
   Constant9_0_impl_instance: Constant_float_8_23_n268_div_65536_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Y => Constant9_0_impl_out);

Delay1No_out_to_Product_0_impl_parent_implementedSystem_port_0_cast <= Delay1No_out;
Delay1No1_out_to_Product_0_impl_parent_implementedSystem_port_1_cast <= Delay1No1_out;
   Product_0_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product_0_impl_out,
                 X => Delay1No_out_to_Product_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No1_out_to_Product_0_impl_parent_implementedSystem_port_1_cast);

SharedReg226_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg226_out;
SharedReg226_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg226_out;
SharedReg226_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg226_out;
SharedReg228_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg228_out;
SharedReg229_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg229_out;
SharedReg229_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg229_out;
SharedReg229_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg229_out;
SharedReg230_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg230_out;
SharedReg231_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg231_out;
SharedReg231_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg231_out;
SharedReg232_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg232_out;
SharedReg232_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg232_out;
SharedReg232_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg232_out;
SharedReg233_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg233_out;
SharedReg233_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg233_out;
SharedReg233_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg233_out;
SharedReg234_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg234_out;
SharedReg234_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg234_out;
SharedReg234_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg234_out;
SharedReg235_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg235_out;
SharedReg235_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg235_out;
SharedReg236_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg236_out;
SharedReg237_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg237_out;
SharedReg237_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg237_out;
SharedReg238_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg238_out;
SharedReg238_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg238_out;
SharedReg239_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg239_out;
SharedReg239_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg239_out;
SharedReg239_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg239_out;
SharedReg240_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg240_out;
SharedReg242_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg242_out;
SharedReg244_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg244_out;
SharedReg244_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg244_out;
SharedReg244_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg244_out;
SharedReg245_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg245_out;
SharedReg245_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg245_out;
SharedReg245_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg245_out;
SharedReg246_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg246_out;
SharedReg246_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg246_out;
SharedReg247_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg247_out;
SharedReg248_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg248_out;
SharedReg248_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg248_out;
SharedReg248_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg248_out;
SharedReg249_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg249_out;
SharedReg249_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg249_out;
SharedReg249_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg249_out;
SharedReg249_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg249_out;
SharedReg250_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg250_out;
SharedReg250_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg250_out;
SharedReg250_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg250_out;
SharedReg251_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg251_out;
SharedReg252_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg252_out;
SharedReg253_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg253_out;
SharedReg254_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg254_out;
SharedReg255_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg255_out;
   MUX_Product_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_55_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg226_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg226_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg232_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg232_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg232_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg233_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg233_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg233_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg234_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg234_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg234_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg235_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg226_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg235_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg236_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg237_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg237_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg238_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg238_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg239_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg239_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg239_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg240_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg228_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg242_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg244_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg244_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg244_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg245_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg245_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg245_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg246_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg246_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg247_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg229_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg248_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg248_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg248_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg249_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg249_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg249_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg249_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg250_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg250_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg250_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg229_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg251_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg252_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg253_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg254_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg255_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_6 => SharedReg229_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg230_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg231_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg231_out_to_MUX_Product_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product_0_impl_0_LUT_out,
                 oMux => MUX_Product_0_impl_0_out);

   Delay1No_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product_0_impl_0_out,
                 Y => Delay1No_out);

SharedReg279_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg279_out;
SharedReg342_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_2_cast <= SharedReg342_out;
SharedReg275_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg275_out;
SharedReg296_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg296_out;
SharedReg317_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg317_out;
SharedReg277_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg277_out;
SharedReg286_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg286_out;
SharedReg278_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg278_out;
SharedReg280_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg280_out;
SharedReg301_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg301_out;
SharedReg285_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg285_out;
SharedReg286_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg286_out;
SharedReg307_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg307_out;
SharedReg284_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg284_out;
SharedReg305_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg305_out;
SharedReg326_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg326_out;
SharedReg279_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg279_out;
SharedReg300_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg300_out;
SharedReg321_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg321_out;
SharedReg283_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg283_out;
SharedReg284_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg284_out;
SharedReg305_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg305_out;
SharedReg326_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg326_out;
SharedReg287_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg287_out;
SharedReg308_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg308_out;
SharedReg329_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg329_out;
SharedReg289_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg289_out;
SharedReg310_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg310_out;
SharedReg331_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg331_out;
SharedReg352_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg352_out;
SharedReg292_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg292_out;
SharedReg290_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg290_out;
SharedReg289_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg289_out;
SharedReg310_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg310_out;
SharedReg288_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg288_out;
SharedReg291_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg291_out;
SharedReg312_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg312_out;
SharedReg354_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg354_out;
SharedReg282_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg282_out;
SharedReg295_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg295_out;
SharedReg316_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg316_out;
SharedReg337_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg337_out;
SharedReg293_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg293_out;
SharedReg314_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg314_out;
SharedReg335_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg335_out;
SharedReg278_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg278_out;
SharedReg299_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg299_out;
SharedReg320_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg320_out;
SharedReg280_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg280_out;
SharedReg281_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg281_out;
SharedReg276_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg276_out;
SharedReg297_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg297_out;
SharedReg339_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg339_out;
SharedReg276_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg276_out;
SharedReg297_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg297_out;
   MUX_Product_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_55_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg279_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg342_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg285_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg286_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg307_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg284_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg305_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg326_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg279_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg300_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg321_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg283_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg275_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg284_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg305_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg326_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg287_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg308_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg329_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg289_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg310_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg331_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg352_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg296_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg292_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg290_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg289_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg310_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg288_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg291_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg312_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg354_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg282_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg295_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg317_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg316_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg337_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg293_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg314_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg335_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg278_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg299_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg320_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg280_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg281_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg277_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg276_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg297_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg339_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg276_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg297_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_6 => SharedReg286_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg278_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg280_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg301_out_to_MUX_Product_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product_0_impl_1_LUT_out,
                 oMux => MUX_Product_0_impl_1_out);

   Delay1No1_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product_0_impl_1_out,
                 Y => Delay1No1_out);

Delay1No2_out_to_Product_2_impl_parent_implementedSystem_port_0_cast <= Delay1No2_out;
Delay1No3_out_to_Product_2_impl_parent_implementedSystem_port_1_cast <= Delay1No3_out;
   Product_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product_2_impl_out,
                 X => Delay1No2_out_to_Product_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No3_out_to_Product_2_impl_parent_implementedSystem_port_1_cast);

SharedReg226_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg226_out;
SharedReg227_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg227_out;
SharedReg227_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg227_out;
SharedReg227_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg227_out;
SharedReg228_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg228_out;
SharedReg228_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg228_out;
SharedReg230_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg230_out;
SharedReg230_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg230_out;
SharedReg231_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg231_out;
SharedReg232_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg232_out;
SharedReg235_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg235_out;
SharedReg235_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg235_out;
SharedReg236_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg236_out;
SharedReg236_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg236_out;
SharedReg237_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg237_out;
SharedReg238_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg238_out;
SharedReg238_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg238_out;
SharedReg239_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg239_out;
SharedReg241_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg241_out;
SharedReg241_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg241_out;
SharedReg241_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg241_out;
SharedReg242_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg242_out;
SharedReg242_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg242_out;
SharedReg242_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg242_out;
SharedReg243_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg243_out;
SharedReg243_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg243_out;
SharedReg243_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg243_out;
SharedReg244_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg244_out;
SharedReg246_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg246_out;
SharedReg247_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg247_out;
SharedReg248_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg248_out;
SharedReg250_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg250_out;
SharedReg251_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg251_out;
SharedReg251_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg251_out;
SharedReg252_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg252_out;
SharedReg252_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg252_out;
SharedReg253_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg253_out;
SharedReg254_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg254_out;
SharedReg254_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg254_out;
SharedReg254_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg254_out;
SharedReg255_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg255_out;
   MUX_Product_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_41_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg226_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg227_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg235_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg235_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg236_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg236_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg237_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg238_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg238_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg239_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg241_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg241_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg227_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg241_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg242_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg242_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg242_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg243_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg243_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg243_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg244_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg246_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg247_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg227_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg248_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg250_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg251_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg251_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg252_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg252_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg253_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg254_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg254_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg254_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg228_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg255_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_5 => SharedReg228_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg230_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg230_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg231_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg232_out_to_MUX_Product_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product_2_impl_0_LUT_out,
                 oMux => MUX_Product_2_impl_0_out);

   Delay1No2_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product_2_impl_0_out,
                 Y => Delay1No2_out);

SharedReg353_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg353_out;
SharedReg300_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg300_out;
SharedReg338_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg338_out;
SharedReg298_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg298_out;
SharedReg340_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg340_out;
SharedReg307_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg307_out;
SharedReg349_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg349_out;
SharedReg299_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg299_out;
SharedReg320_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg320_out;
SharedReg341_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg341_out;
SharedReg322_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg322_out;
SharedReg306_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg306_out;
SharedReg327_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg327_out;
SharedReg328_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg328_out;
SharedReg347_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg347_out;
SharedReg342_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg342_out;
SharedReg304_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg304_out;
SharedReg294_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg294_out;
SharedReg315_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg315_out;
SharedReg336_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg336_out;
SharedReg311_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg311_out;
SharedReg332_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg332_out;
SharedReg331_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg331_out;
SharedReg352_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg352_out;
SharedReg309_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg309_out;
SharedReg333_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg333_out;
Delay123No_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_27_cast <= Delay123No_out;
Delay123No1_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_28_cast <= Delay123No1_out;
Delay123No2_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_29_cast <= Delay123No2_out;
SharedReg303_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg303_out;
SharedReg324_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg324_out;
SharedReg358_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_32_cast <= SharedReg358_out;
SharedReg301_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg301_out;
SharedReg322_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg322_out;
SharedReg302_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg302_out;
SharedReg318_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg318_out;
SharedReg277_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg277_out;
SharedReg298_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg298_out;
SharedReg340_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg340_out;
SharedReg318_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg318_out;
SharedReg339_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg339_out;
   MUX_Product_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_41_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg353_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg300_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg322_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg306_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg327_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg328_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg347_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg342_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg304_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg294_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg315_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg336_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg338_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg311_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg332_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg331_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg352_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg309_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg333_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => Delay123No_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => Delay123No1_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => Delay123No2_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg303_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg298_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg324_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg358_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg301_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg322_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg302_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg318_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg277_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg298_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg340_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg318_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg340_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg339_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_5 => SharedReg307_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg349_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg299_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg320_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg341_out_to_MUX_Product_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product_2_impl_1_LUT_out,
                 oMux => MUX_Product_2_impl_1_out);

   Delay1No3_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product_2_impl_1_out,
                 Y => Delay1No3_out);

Delay1No4_out_to_Product1_2_impl_parent_implementedSystem_port_0_cast <= Delay1No4_out;
Delay1No5_out_to_Product1_2_impl_parent_implementedSystem_port_1_cast <= Delay1No5_out;
   Product1_2_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product1_2_impl_out,
                 X => Delay1No4_out_to_Product1_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No5_out_to_Product1_2_impl_parent_implementedSystem_port_1_cast);

SharedReg227_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg227_out;
SharedReg229_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg229_out;
SharedReg231_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg231_out;
SharedReg233_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg233_out;
SharedReg234_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg234_out;
SharedReg236_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg236_out;
SharedReg240_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg240_out;
SharedReg240_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg240_out;
SharedReg240_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg240_out;
SharedReg241_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg241_out;
SharedReg245_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg245_out;
SharedReg246_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg246_out;
SharedReg247_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg247_out;
SharedReg251_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg251_out;
SharedReg252_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg252_out;
SharedReg253_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg253_out;
SharedReg253_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg253_out;
SharedReg255_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg255_out;
SharedReg255_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg255_out;
   MUX_Product1_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_19_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg227_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg229_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg245_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg246_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg247_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg251_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg252_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg253_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg253_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg255_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg255_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_2 => SharedReg231_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg233_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg234_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg236_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg240_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg240_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg240_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg241_out_to_MUX_Product1_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product1_2_impl_0_LUT_out,
                 oMux => MUX_Product1_2_impl_0_out);

   Delay1No4_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product1_2_impl_0_out,
                 Y => Delay1No4_out);

SharedReg321_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg321_out;
SharedReg319_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg319_out;
SharedReg328_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg328_out;
SharedReg343_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg343_out;
SharedReg348_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg348_out;
SharedReg325_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg325_out;
SharedReg346_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg346_out;
SharedReg347_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg347_out;
SharedReg350_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg350_out;
SharedReg313_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg313_out;
SharedReg334_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg334_out;
SharedReg355_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg355_out;
SharedReg357_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg357_out;
SharedReg351_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg351_out;
SharedReg356_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg356_out;
SharedReg341_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg341_out;
SharedReg323_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg323_out;
SharedReg344_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg344_out;
SharedReg319_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg319_out;
   MUX_Product1_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_19_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg321_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg319_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg334_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg355_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg357_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg351_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg356_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg341_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg323_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg344_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg319_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_2 => SharedReg328_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg343_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg348_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_5 => SharedReg325_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_6 => SharedReg346_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg347_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg350_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg313_out_to_MUX_Product1_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => MUX_Product1_2_impl_1_LUT_out,
                 oMux => MUX_Product1_2_impl_1_out);

   Delay1No5_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product1_2_impl_1_out,
                 Y => Delay1No5_out);

Delay1No6_out_to_Product10_3_impl_parent_implementedSystem_port_0_cast <= Delay1No6_out;
Delay1No7_out_to_Product10_3_impl_parent_implementedSystem_port_1_cast <= Delay1No7_out;
   Product10_3_impl_instance: FPMultiplier_in_8_23_8_23_out_8_23_mult_X_mult_Y_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Product10_3_impl_out,
                 X => Delay1No6_out_to_Product10_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No7_out_to_Product10_3_impl_parent_implementedSystem_port_1_cast);

SharedReg228_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg228_out;
SharedReg230_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg230_out;
SharedReg237_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg237_out;
SharedReg243_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg243_out;
SharedReg247_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg247_out;
   MUX_Product10_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg228_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg230_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_2 => SharedReg237_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg243_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg247_out_to_MUX_Product10_3_impl_0_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Product10_3_impl_0_LUT_out,
                 oMux => MUX_Product10_3_impl_0_out);

   Delay1No6_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product10_3_impl_0_out,
                 Y => Delay1No6_out);

SharedReg349_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg349_out;
SharedReg330_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg330_out;
Delay123No3_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_3_cast <= Delay123No3_out;
SharedReg345_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg345_out;
SharedReg343_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg343_out;
   MUX_Product10_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_5_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg349_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg330_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_2 => Delay123No3_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_3 => SharedReg345_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_4 => SharedReg343_out_to_MUX_Product10_3_impl_1_parent_implementedSystem_port_5_cast,
                 iSel => MUX_Product10_3_impl_1_LUT_out,
                 oMux => MUX_Product10_3_impl_1_out);

   Delay1No7_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Product10_3_impl_1_out,
                 Y => Delay1No7_out);

Delay1No8_out_to_Sum10_0_impl_parent_implementedSystem_port_0_cast <= Delay1No8_out;
Delay1No9_out_to_Sum10_0_impl_parent_implementedSystem_port_1_cast <= Delay1No9_out;
   Sum10_0_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Sum10_0_impl_out,
                 X => Delay1No8_out_to_Sum10_0_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No9_out_to_Sum10_0_impl_parent_implementedSystem_port_1_cast);

SharedReg170_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_1_cast <= SharedReg170_out;
SharedReg_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_2_cast <= SharedReg_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_3_cast <= SharedReg275_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_4_cast <= SharedReg275_out;
SharedReg191_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_5_cast <= SharedReg191_out;
SharedReg114_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_6_cast <= SharedReg114_out;
SharedReg59_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_7_cast <= SharedReg59_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_8_cast <= SharedReg275_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_9_cast <= SharedReg275_out;
SharedReg118_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_10_cast <= SharedReg118_out;
SharedReg80_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_11_cast <= SharedReg80_out;
SharedReg256_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_12_cast <= SharedReg256_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_13_cast <= SharedReg275_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_14_cast <= SharedReg275_out;
SharedReg133_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_15_cast <= SharedReg133_out;
SharedReg4_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_16_cast <= SharedReg4_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_17_cast <= SharedReg275_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_18_cast <= SharedReg275_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_19_cast <= SharedReg275_out;
SharedReg25_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_20_cast <= SharedReg25_out;
SharedReg174_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_21_cast <= SharedReg174_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_22_cast <= SharedReg275_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_23_cast <= SharedReg275_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_24_cast <= SharedReg275_out;
SharedReg63_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_25_cast <= SharedReg63_out;
SharedReg23_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_26_cast <= SharedReg23_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_27_cast <= SharedReg275_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_28_cast <= SharedReg275_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_29_cast <= SharedReg275_out;
SharedReg178_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_30_cast <= SharedReg178_out;
SharedReg185_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_31_cast <= SharedReg185_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_32_cast <= SharedReg275_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_33_cast <= SharedReg275_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_34_cast <= SharedReg275_out;
SharedReg8_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_35_cast <= SharedReg8_out;
SharedReg122_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_36_cast <= SharedReg122_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_37_cast <= SharedReg275_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_38_cast <= SharedReg275_out;
SharedReg19_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_39_cast <= SharedReg19_out;
SharedReg73_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_40_cast <= SharedReg73_out;
SharedReg79_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_41_cast <= SharedReg79_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_42_cast <= SharedReg275_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_43_cast <= SharedReg275_out;
SharedReg126_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_44_cast <= SharedReg126_out;
SharedReg197_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_45_cast <= SharedReg197_out;
SharedReg16_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_46_cast <= SharedReg16_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_47_cast <= SharedReg275_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_48_cast <= SharedReg275_out;
SharedReg190_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_49_cast <= SharedReg190_out;
SharedReg67_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_50_cast <= SharedReg67_out;
SharedReg12_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_51_cast <= SharedReg12_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_52_cast <= SharedReg275_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_53_cast <= SharedReg275_out;
SharedReg139_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_54_cast <= SharedReg139_out;
SharedReg71_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_55_cast <= SharedReg71_out;
SharedReg182_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_56_cast <= SharedReg182_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_57_cast <= SharedReg275_out;
SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_58_cast <= SharedReg275_out;
SharedReg131_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_59_cast <= SharedReg131_out;
   MUX_Sum10_0_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg170_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg80_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg256_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg133_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg4_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg25_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg174_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg63_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg23_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg178_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg185_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg8_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg122_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg19_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg73_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg191_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg79_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg126_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg197_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg16_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg190_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg67_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg114_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg12_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg139_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg71_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg182_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg131_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_59_cast,
                 iS_6 => SharedReg59_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg275_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg118_out_to_MUX_Sum10_0_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum10_0_impl_0_out);

   Delay1No8_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum10_0_impl_0_out,
                 Y => Delay1No8_out);

SharedReg168_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_1_cast <= SharedReg168_out;
Delay871No1_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_2_cast <= Delay871No1_out;
SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_3_cast <= SharedReg256_out;
SharedReg260_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_4_cast <= SharedReg260_out;
SharedReg144_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_5_cast <= SharedReg144_out;
SharedReg224_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_6_cast <= SharedReg224_out;
SharedReg53_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_7_cast <= SharedReg53_out;
SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_8_cast <= SharedReg256_out;
SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_9_cast <= SharedReg256_out;
SharedReg220_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_10_cast <= SharedReg220_out;
SharedReg29_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_11_cast <= SharedReg29_out;
SharedReg264_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_12_cast <= SharedReg264_out;
SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_13_cast <= SharedReg256_out;
SharedReg267_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_14_cast <= SharedReg267_out;
SharedReg204_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_15_cast <= SharedReg204_out;
SharedReg108_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_16_cast <= SharedReg108_out;
SharedReg257_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_17_cast <= SharedReg257_out;
SharedReg259_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_18_cast <= SharedReg259_out;
SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_19_cast <= SharedReg256_out;
SharedReg84_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_20_cast <= SharedReg84_out;
SharedReg164_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_21_cast <= SharedReg164_out;
SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_22_cast <= SharedReg256_out;
SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_23_cast <= SharedReg256_out;
SharedReg264_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_24_cast <= SharedReg264_out;
SharedReg50_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_25_cast <= SharedReg50_out;
SharedReg89_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_26_cast <= SharedReg89_out;
SharedReg258_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_27_cast <= SharedReg258_out;
SharedReg262_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_28_cast <= SharedReg262_out;
SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_29_cast <= SharedReg256_out;
SharedReg160_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_30_cast <= SharedReg160_out;
SharedReg152_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_31_cast <= SharedReg152_out;
SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_32_cast <= SharedReg256_out;
SharedReg263_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_33_cast <= SharedReg263_out;
SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_34_cast <= SharedReg256_out;
SharedReg105_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_35_cast <= SharedReg105_out;
SharedReg217_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_36_cast <= SharedReg217_out;
SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_37_cast <= SharedReg256_out;
SharedReg261_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_38_cast <= SharedReg261_out;
SharedReg93_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_39_cast <= SharedReg93_out;
SharedReg38_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_40_cast <= SharedReg38_out;
SharedReg35_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_41_cast <= SharedReg35_out;
SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_42_cast <= SharedReg256_out;
SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_43_cast <= SharedReg256_out;
SharedReg213_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_44_cast <= SharedReg213_out;
SharedReg143_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_45_cast <= SharedReg143_out;
SharedReg97_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_46_cast <= SharedReg97_out;
SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_47_cast <= SharedReg256_out;
SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_48_cast <= SharedReg256_out;
SharedReg149_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_49_cast <= SharedReg149_out;
SharedReg46_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_50_cast <= SharedReg46_out;
SharedReg101_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_51_cast <= SharedReg101_out;
SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_52_cast <= SharedReg256_out;
SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_53_cast <= SharedReg256_out;
SharedReg202_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_54_cast <= SharedReg202_out;
SharedReg42_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_55_cast <= SharedReg42_out;
SharedReg157_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_56_cast <= SharedReg157_out;
SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_57_cast <= SharedReg256_out;
SharedReg260_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_58_cast <= SharedReg260_out;
SharedReg210_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_59_cast <= SharedReg210_out;
   MUX_Sum10_0_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg168_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => Delay871No1_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg29_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg264_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg267_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg204_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg108_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg257_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg259_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg84_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg164_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg264_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg50_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg89_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg258_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg262_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg160_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg260_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg152_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg263_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg105_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg217_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg261_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg93_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg38_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg144_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg35_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg213_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg143_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg97_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg149_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg46_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg224_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg101_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg202_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg42_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg157_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg260_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg210_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_59_cast,
                 iS_6 => SharedReg53_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg256_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg220_out_to_MUX_Sum10_0_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum10_0_impl_1_out);

   Delay1No9_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum10_0_impl_1_out,
                 Y => Delay1No9_out);

Delay1No10_out_to_Sum10_1_impl_parent_implementedSystem_port_0_cast <= Delay1No10_out;
Delay1No11_out_to_Sum10_1_impl_parent_implementedSystem_port_1_cast <= Delay1No11_out;
   Sum10_1_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Sum10_1_impl_out,
                 X => Delay1No10_out_to_Sum10_1_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No11_out_to_Sum10_1_impl_parent_implementedSystem_port_1_cast);

SharedReg27_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_1_cast <= SharedReg27_out;
SharedReg72_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_2_cast <= SharedReg72_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_3_cast <= SharedReg296_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_4_cast <= SharedReg296_out;
SharedReg21_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_5_cast <= SharedReg21_out;
SharedReg123_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_6_cast <= SharedReg123_out;
SharedReg68_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_7_cast <= SharedReg68_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_8_cast <= SharedReg296_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_9_cast <= SharedReg296_out;
SharedReg196_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_10_cast <= SharedReg196_out;
SharedReg127_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_11_cast <= SharedReg127_out;
SharedReg13_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_12_cast <= SharedReg13_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_13_cast <= SharedReg296_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_14_cast <= SharedReg296_out;
SharedReg187_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_15_cast <= SharedReg187_out;
SharedReg1_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_16_cast <= SharedReg1_out;
SharedReg56_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_17_cast <= SharedReg56_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_18_cast <= SharedReg296_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_19_cast <= SharedReg296_out;
SharedReg22_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_20_cast <= SharedReg22_out;
SharedReg171_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_21_cast <= SharedReg171_out;
SharedReg115_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_22_cast <= SharedReg115_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_23_cast <= SharedReg296_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_24_cast <= SharedReg296_out;
SharedReg175_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_25_cast <= SharedReg175_out;
SharedReg137_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_26_cast <= SharedReg137_out;
SharedReg256_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_27_cast <= SharedReg256_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_28_cast <= SharedReg296_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_29_cast <= SharedReg296_out;
SharedReg189_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_30_cast <= SharedReg189_out;
SharedReg60_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_31_cast <= SharedReg60_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_32_cast <= SharedReg296_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_33_cast <= SharedReg296_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_34_cast <= SharedReg296_out;
SharedReg81_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_35_cast <= SharedReg81_out;
SharedReg5_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_36_cast <= SharedReg5_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_37_cast <= SharedReg296_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_38_cast <= SharedReg296_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_39_cast <= SharedReg296_out;
SharedReg119_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_40_cast <= SharedReg119_out;
SharedReg79_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_41_cast <= SharedReg79_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_42_cast <= SharedReg296_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_43_cast <= SharedReg296_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_44_cast <= SharedReg296_out;
SharedReg9_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_45_cast <= SharedReg9_out;
SharedReg16_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_46_cast <= SharedReg16_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_47_cast <= SharedReg296_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_48_cast <= SharedReg296_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_49_cast <= SharedReg296_out;
SharedReg64_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_50_cast <= SharedReg64_out;
SharedReg179_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_51_cast <= SharedReg179_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_52_cast <= SharedReg296_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_53_cast <= SharedReg296_out;
SharedReg75_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_54_cast <= SharedReg75_out;
SharedReg130_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_55_cast <= SharedReg130_out;
SharedReg136_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_56_cast <= SharedReg136_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_57_cast <= SharedReg296_out;
SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_58_cast <= SharedReg296_out;
SharedReg183_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_59_cast <= SharedReg183_out;
   MUX_Sum10_1_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg27_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg72_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg127_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg13_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg187_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg1_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg56_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg22_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg171_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg115_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg175_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg137_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg256_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg189_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg60_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg81_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg5_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg119_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg21_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg79_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg9_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg16_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg64_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg123_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg179_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg75_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg130_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg136_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg183_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_59_cast,
                 iS_6 => SharedReg68_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg296_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg196_out_to_MUX_Sum10_1_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum10_1_impl_0_out);

   Delay1No10_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum10_1_impl_0_out,
                 Y => Delay1No10_out);

SharedReg200_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_1_cast <= SharedReg200_out;
SharedReg154_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_2_cast <= SharedReg154_out;
SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_3_cast <= SharedReg264_out;
SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_4_cast <= SharedReg256_out;
SharedReg206_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_5_cast <= SharedReg206_out;
SharedReg102_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_6_cast <= SharedReg102_out;
SharedReg158_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_7_cast <= SharedReg158_out;
SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_8_cast <= SharedReg264_out;
SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_9_cast <= SharedReg264_out;
SharedReg32_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_10_cast <= SharedReg32_out;
SharedReg98_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_11_cast <= SharedReg98_out;
SharedReg214_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_12_cast <= SharedReg214_out;
SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_13_cast <= SharedReg264_out;
SharedReg260_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_14_cast <= SharedReg260_out;
SharedReg40_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_15_cast <= SharedReg40_out;
SharedReg225_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_16_cast <= SharedReg225_out;
Delay871No2_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_17_cast <= Delay871No2_out;
SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_18_cast <= SharedReg256_out;
SharedReg260_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_19_cast <= SharedReg260_out;
SharedReg201_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_20_cast <= SharedReg201_out;
SharedReg54_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_21_cast <= SharedReg54_out;
SharedReg109_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_22_cast <= SharedReg109_out;
SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_23_cast <= SharedReg264_out;
SharedReg271_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_24_cast <= SharedReg271_out;
SharedReg50_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_25_cast <= SharedReg50_out;
SharedReg85_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_26_cast <= SharedReg85_out;
SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_27_cast <= SharedReg264_out;
SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_28_cast <= SharedReg256_out;
SharedReg267_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_29_cast <= SharedReg267_out;
SharedReg34_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_30_cast <= SharedReg34_out;
SharedReg165_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_31_cast <= SharedReg165_out;
SharedReg257_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_32_cast <= SharedReg257_out;
SharedReg268_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_33_cast <= SharedReg268_out;
SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_34_cast <= SharedReg264_out;
SharedReg141_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_35_cast <= SharedReg141_out;
SharedReg221_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_36_cast <= SharedReg221_out;
SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_37_cast <= SharedReg264_out;
SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_38_cast <= SharedReg256_out;
SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_39_cast <= SharedReg264_out;
SharedReg106_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_40_cast <= SharedReg106_out;
SharedReg146_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_41_cast <= SharedReg146_out;
SharedReg258_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_42_cast <= SharedReg258_out;
SharedReg262_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_43_cast <= SharedReg262_out;
SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_44_cast <= SharedReg256_out;
SharedReg218_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_45_cast <= SharedReg218_out;
SharedReg209_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_46_cast <= SharedReg209_out;
SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_47_cast <= SharedReg264_out;
SharedReg263_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_48_cast <= SharedReg263_out;
SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_49_cast <= SharedReg256_out;
SharedReg161_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_50_cast <= SharedReg161_out;
SharedReg47_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_51_cast <= SharedReg47_out;
SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_52_cast <= SharedReg264_out;
SharedReg261_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_53_cast <= SharedReg261_out;
SharedReg150_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_54_cast <= SharedReg150_out;
SharedReg94_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_55_cast <= SharedReg94_out;
SharedReg91_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_56_cast <= SharedReg91_out;
SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_57_cast <= SharedReg264_out;
SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_58_cast <= SharedReg256_out;
SharedReg43_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_59_cast <= SharedReg43_out;
   MUX_Sum10_1_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg200_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg154_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg98_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg214_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg260_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg40_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg225_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => Delay871No2_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg260_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg201_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg54_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg109_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg271_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg50_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg85_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg267_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg34_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg165_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg257_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg268_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg141_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg221_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg106_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg206_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg146_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg258_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg262_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg218_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg209_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg263_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg161_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg102_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg47_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg261_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg150_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg94_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg91_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg256_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg43_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_59_cast,
                 iS_6 => SharedReg158_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg264_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg32_out_to_MUX_Sum10_1_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum10_1_impl_1_out);

   Delay1No11_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum10_1_impl_1_out,
                 Y => Delay1No11_out);

Delay1No12_out_to_Sum10_2_impl_parent_implementedSystem_port_0_cast <= Delay1No12_out;
Delay1No13_out_to_Sum10_2_impl_parent_implementedSystem_port_1_cast <= Delay1No13_out;
   Sum10_2_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Sum10_2_impl_out,
                 X => Delay1No12_out_to_Sum10_2_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No13_out_to_Sum10_2_impl_parent_implementedSystem_port_1_cast);

SharedReg65_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_1_cast <= SharedReg65_out;
SharedReg72_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_2_cast <= SharedReg72_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_3_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_4_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_5_cast <= SharedReg317_out;
SharedReg120_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_6_cast <= SharedReg120_out;
SharedReg10_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_7_cast <= SharedReg10_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_8_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_9_cast <= SharedReg317_out;
SharedReg132_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_10_cast <= SharedReg132_out;
SharedReg186_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_11_cast <= SharedReg186_out;
SharedReg193_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_12_cast <= SharedReg193_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_13_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_14_cast <= SharedReg317_out;
SharedReg14_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_15_cast <= SharedReg14_out;
SharedReg83_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_16_cast <= SharedReg83_out;
SharedReg129_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_17_cast <= SharedReg129_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_18_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_19_cast <= SharedReg317_out;
SharedReg77_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_20_cast <= SharedReg77_out;
SharedReg180_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_21_cast <= SharedReg180_out;
SharedReg124_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_22_cast <= SharedReg124_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_23_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_24_cast <= SharedReg317_out;
SharedReg26_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_25_cast <= SharedReg26_out;
SharedReg184_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_26_cast <= SharedReg184_out;
SharedReg69_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_27_cast <= SharedReg69_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_28_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_29_cast <= SharedReg317_out;
SharedReg18_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_30_cast <= SharedReg18_out;
SharedReg57_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_31_cast <= SharedReg57_out;
SharedReg112_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_32_cast <= SharedReg112_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_33_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_34_cast <= SharedReg317_out;
SharedReg78_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_35_cast <= SharedReg78_out;
SharedReg2_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_36_cast <= SharedReg2_out;
SharedReg172_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_37_cast <= SharedReg172_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_38_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_39_cast <= SharedReg317_out;
SharedReg6_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_40_cast <= SharedReg6_out;
SharedReg194_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_41_cast <= SharedReg194_out;
SharedReg264_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_42_cast <= SharedReg264_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_43_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_44_cast <= SharedReg317_out;
SharedReg20_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_45_cast <= SharedReg20_out;
SharedReg116_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_46_cast <= SharedReg116_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_47_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_48_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_49_cast <= SharedReg317_out;
SharedReg138_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_50_cast <= SharedReg138_out;
SharedReg61_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_51_cast <= SharedReg61_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_52_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_53_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_54_cast <= SharedReg317_out;
SharedReg176_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_55_cast <= SharedReg176_out;
SharedReg136_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_56_cast <= SharedReg136_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_57_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_58_cast <= SharedReg317_out;
SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_59_cast <= SharedReg317_out;
   MUX_Sum10_2_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg65_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg72_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg186_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg193_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg14_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg83_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg129_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg77_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg180_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg124_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg26_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg184_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg69_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg18_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg57_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg112_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg78_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg2_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg172_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg6_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg194_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg264_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg20_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg116_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg138_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg120_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg61_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg176_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg136_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_59_cast,
                 iS_6 => SharedReg10_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg317_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg132_out_to_MUX_Sum10_2_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum10_2_impl_0_out);

   Delay1No12_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum10_2_impl_0_out,
                 Y => Delay1No12_out);

SharedReg48_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_1_cast <= SharedReg48_out;
SharedReg39_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_2_cast <= SharedReg39_out;
SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_3_cast <= SharedReg271_out;
SharedReg263_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_4_cast <= SharedReg263_out;
SharedReg256_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_5_cast <= SharedReg256_out;
SharedReg219_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_6_cast <= SharedReg219_out;
SharedReg103_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_7_cast <= SharedReg103_out;
SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_8_cast <= SharedReg271_out;
SharedReg261_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_9_cast <= SharedReg261_out;
SharedReg207_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_10_cast <= SharedReg207_out;
SharedReg151_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_11_cast <= SharedReg151_out;
SharedReg148_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_12_cast <= SharedReg148_out;
SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_13_cast <= SharedReg271_out;
SharedReg256_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_14_cast <= SharedReg256_out;
SharedReg99_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_15_cast <= SharedReg99_out;
SharedReg30_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_16_cast <= SharedReg30_out;
SharedReg211_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_17_cast <= SharedReg211_out;
SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_18_cast <= SharedReg264_out;
SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_19_cast <= SharedReg264_out;
SharedReg36_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_20_cast <= SharedReg36_out;
SharedReg159_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_21_cast <= SharedReg159_out;
SharedReg215_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_22_cast <= SharedReg215_out;
SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_23_cast <= SharedReg271_out;
SharedReg274_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_24_cast <= SharedReg274_out;
SharedReg88_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_25_cast <= SharedReg88_out;
SharedReg155_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_26_cast <= SharedReg155_out;
SharedReg44_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_27_cast <= SharedReg44_out;
SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_28_cast <= SharedReg264_out;
SharedReg269_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_29_cast <= SharedReg269_out;
SharedReg96_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_30_cast <= SharedReg96_out;
SharedReg55_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_31_cast <= SharedReg55_out;
Delay872No_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_32_cast <= Delay872No_out;
SharedReg256_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_33_cast <= SharedReg256_out;
SharedReg260_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_34_cast <= SharedReg260_out;
SharedReg31_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_35_cast <= SharedReg31_out;
SharedReg110_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_36_cast <= SharedReg110_out;
SharedReg166_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_37_cast <= SharedReg166_out;
SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_38_cast <= SharedReg264_out;
SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_39_cast <= SharedReg271_out;
SharedReg106_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_40_cast <= SharedReg106_out;
SharedReg142_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_41_cast <= SharedReg142_out;
SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_42_cast <= SharedReg271_out;
SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_43_cast <= SharedReg264_out;
SharedReg267_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_44_cast <= SharedReg267_out;
SharedReg90_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_45_cast <= SharedReg90_out;
SharedReg222_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_46_cast <= SharedReg222_out;
SharedReg265_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_47_cast <= SharedReg265_out;
SharedReg268_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_48_cast <= SharedReg268_out;
SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_49_cast <= SharedReg264_out;
SharedReg198_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_50_cast <= SharedReg198_out;
SharedReg51_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_51_cast <= SharedReg51_out;
SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_52_cast <= SharedReg271_out;
SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_53_cast <= SharedReg264_out;
SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_54_cast <= SharedReg264_out;
SharedReg163_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_55_cast <= SharedReg163_out;
SharedReg203_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_56_cast <= SharedReg203_out;
SharedReg258_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_57_cast <= SharedReg258_out;
SharedReg262_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_58_cast <= SharedReg262_out;
SharedReg256_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_59_cast <= SharedReg256_out;
   MUX_Sum10_2_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg48_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg39_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg151_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg148_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg256_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg99_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg30_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg211_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg36_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg159_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg215_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg274_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg88_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg155_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg44_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg269_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg96_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg263_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg55_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => Delay872No_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg256_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg260_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg31_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg110_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg166_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg106_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg256_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg142_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg267_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg90_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg222_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg265_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg268_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg198_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg219_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg51_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg264_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg163_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg203_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg258_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg262_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg256_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_59_cast,
                 iS_6 => SharedReg103_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg271_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg261_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg207_out_to_MUX_Sum10_2_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum10_2_impl_1_out);

   Delay1No13_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum10_2_impl_1_out,
                 Y => Delay1No13_out);

Delay1No14_out_to_Sum10_3_impl_parent_implementedSystem_port_0_cast <= Delay1No14_out;
Delay1No15_out_to_Sum10_3_impl_parent_implementedSystem_port_1_cast <= Delay1No15_out;
   Sum10_3_impl_instance: FPGenericAddSub_wE_8_wF_23_subX_false_subY_false_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Sum10_3_impl_out,
                 X => Delay1No14_out_to_Sum10_3_impl_parent_implementedSystem_port_0_cast,
                 Y => Delay1No15_out_to_Sum10_3_impl_parent_implementedSystem_port_1_cast);

SharedReg173_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_1_cast <= SharedReg173_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_2_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_3_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_4_cast <= SharedReg338_out;
SharedReg195_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_5_cast <= SharedReg195_out;
SharedReg117_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_6_cast <= SharedReg117_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_7_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_8_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_9_cast <= SharedReg338_out;
SharedReg7_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_10_cast <= SharedReg7_out;
SharedReg192_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_11_cast <= SharedReg192_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_12_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_13_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_14_cast <= SharedReg338_out;
SharedReg121_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_15_cast <= SharedReg121_out;
SharedReg128_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_16_cast <= SharedReg128_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_17_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_18_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_19_cast <= SharedReg338_out;
SharedReg177_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_20_cast <= SharedReg177_out;
SharedReg66_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_21_cast <= SharedReg66_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_22_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_23_cast <= SharedReg338_out;
SharedReg188_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_24_cast <= SharedReg188_out;
SharedReg17_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_25_cast <= SharedReg17_out;
SharedReg23_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_26_cast <= SharedReg23_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_27_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_28_cast <= SharedReg338_out;
SharedReg70_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_29_cast <= SharedReg70_out;
SharedReg140_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_30_cast <= SharedReg140_out;
SharedReg185_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_31_cast <= SharedReg185_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_32_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_33_cast <= SharedReg338_out;
SharedReg134_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_34_cast <= SharedReg134_out;
SharedReg11_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_35_cast <= SharedReg11_out;
SharedReg181_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_36_cast <= SharedReg181_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_37_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_38_cast <= SharedReg338_out;
SharedReg82_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_39_cast <= SharedReg82_out;
SharedReg15_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_40_cast <= SharedReg15_out;
SharedReg125_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_41_cast <= SharedReg125_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_42_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_43_cast <= SharedReg338_out;
SharedReg74_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_44_cast <= SharedReg74_out;
SharedReg113_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_45_cast <= SharedReg113_out;
SharedReg169_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_46_cast <= SharedReg169_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_47_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_48_cast <= SharedReg338_out;
SharedReg135_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_49_cast <= SharedReg135_out;
SharedReg58_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_50_cast <= SharedReg58_out;
SharedReg3_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_51_cast <= SharedReg3_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_52_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_53_cast <= SharedReg338_out;
SharedReg62_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_54_cast <= SharedReg62_out;
SharedReg24_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_55_cast <= SharedReg24_out;
SharedReg256_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_56_cast <= SharedReg256_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_57_cast <= SharedReg338_out;
SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_58_cast <= SharedReg338_out;
SharedReg76_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_59_cast <= SharedReg76_out;
   MUX_Sum10_3_impl_0_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg173_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg192_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg121_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg128_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_17_cast,
                 iS_17 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg177_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg66_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_22_cast,
                 iS_22 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg188_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg17_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg23_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg70_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg140_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg185_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg134_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg11_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg181_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg82_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg15_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg195_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg125_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg74_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg113_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_45_cast,
                 iS_45 => SharedReg169_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg135_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg58_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg117_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg3_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg62_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg24_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg256_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg76_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_59_cast,
                 iS_6 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg338_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg7_out_to_MUX_Sum10_3_impl_0_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum10_3_impl_0_out);

   Delay1No14_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum10_3_impl_0_out,
                 Y => Delay1No14_out);

SharedReg52_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_1_cast <= SharedReg52_out;
SharedReg265_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_2_cast <= SharedReg265_out;
SharedReg273_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_3_cast <= SharedReg273_out;
SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_4_cast <= SharedReg264_out;
SharedReg28_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_5_cast <= SharedReg28_out;
SharedReg107_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_6_cast <= SharedReg107_out;
SharedReg256_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_7_cast <= SharedReg256_out;
SharedReg274_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_8_cast <= SharedReg274_out;
SharedReg274_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_9_cast <= SharedReg274_out;
SharedReg220_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_10_cast <= SharedReg220_out;
SharedReg33_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_11_cast <= SharedReg33_out;
SharedReg266_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_12_cast <= SharedReg266_out;
SharedReg270_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_13_cast <= SharedReg270_out;
SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_14_cast <= SharedReg264_out;
SharedReg104_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_15_cast <= SharedReg104_out;
SharedReg95_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_16_cast <= SharedReg95_out;
SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_17_cast <= SharedReg264_out;
Delay47No7_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_18_cast <= Delay47No7_out;
SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_19_cast <= SharedReg271_out;
SharedReg49_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_20_cast <= SharedReg49_out;
SharedReg159_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_21_cast <= SharedReg159_out;
SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_22_cast <= SharedReg264_out;
Delay15No6_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_23_cast <= Delay15No6_out;
SharedReg37_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_24_cast <= SharedReg37_out;
SharedReg208_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_25_cast <= SharedReg208_out;
SharedReg205_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_26_cast <= SharedReg205_out;
SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_27_cast <= SharedReg271_out;
SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_28_cast <= SharedReg271_out;
SharedReg156_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_29_cast <= SharedReg156_out;
SharedReg86_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_30_cast <= SharedReg86_out;
SharedReg41_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_31_cast <= SharedReg41_out;
SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_32_cast <= SharedReg264_out;
SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_33_cast <= SharedReg264_out;
SharedReg92_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_34_cast <= SharedReg92_out;
SharedReg216_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_35_cast <= SharedReg216_out;
SharedReg45_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_36_cast <= SharedReg45_out;
SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_37_cast <= SharedReg271_out;
SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_38_cast <= SharedReg271_out;
SharedReg145_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_39_cast <= SharedReg145_out;
SharedReg212_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_40_cast <= SharedReg212_out;
SharedReg100_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_41_cast <= SharedReg100_out;
SharedReg274_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_42_cast <= SharedReg274_out;
SharedReg260_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_43_cast <= SharedReg260_out;
SharedReg153_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_44_cast <= SharedReg153_out;
SharedReg111_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_45_cast <= SharedReg111_out;
Delay871No_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_46_cast <= Delay871No_out;
SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_47_cast <= SharedReg271_out;
SharedReg260_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_48_cast <= SharedReg260_out;
SharedReg87_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_49_cast <= SharedReg87_out;
SharedReg167_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_50_cast <= SharedReg167_out;
SharedReg223_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_51_cast <= SharedReg223_out;
SharedReg274_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_52_cast <= SharedReg274_out;
SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_53_cast <= SharedReg271_out;
SharedReg162_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_54_cast <= SharedReg162_out;
SharedReg199_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_55_cast <= SharedReg199_out;
SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_56_cast <= SharedReg264_out;
SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_57_cast <= SharedReg271_out;
SharedReg272_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_58_cast <= SharedReg272_out;
SharedReg147_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_59_cast <= SharedReg147_out;
   MUX_Sum10_3_impl_1_instance: Mux_sign_1_wordsize_34_numberOfInputs_59_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 iS_0 => SharedReg52_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_1_cast,
                 iS_1 => SharedReg265_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_2_cast,
                 iS_10 => SharedReg33_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_11_cast,
                 iS_11 => SharedReg266_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_12_cast,
                 iS_12 => SharedReg270_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_13_cast,
                 iS_13 => SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_14_cast,
                 iS_14 => SharedReg104_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_15_cast,
                 iS_15 => SharedReg95_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_16_cast,
                 iS_16 => SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_17_cast,
                 iS_17 => Delay47No7_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_18_cast,
                 iS_18 => SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_19_cast,
                 iS_19 => SharedReg49_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_20_cast,
                 iS_2 => SharedReg273_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_3_cast,
                 iS_20 => SharedReg159_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_21_cast,
                 iS_21 => SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_22_cast,
                 iS_22 => Delay15No6_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_23_cast,
                 iS_23 => SharedReg37_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_24_cast,
                 iS_24 => SharedReg208_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_25_cast,
                 iS_25 => SharedReg205_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_26_cast,
                 iS_26 => SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_27_cast,
                 iS_27 => SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_28_cast,
                 iS_28 => SharedReg156_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_29_cast,
                 iS_29 => SharedReg86_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_30_cast,
                 iS_3 => SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_4_cast,
                 iS_30 => SharedReg41_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_31_cast,
                 iS_31 => SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_32_cast,
                 iS_32 => SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_33_cast,
                 iS_33 => SharedReg92_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_34_cast,
                 iS_34 => SharedReg216_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_35_cast,
                 iS_35 => SharedReg45_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_36_cast,
                 iS_36 => SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_37_cast,
                 iS_37 => SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_38_cast,
                 iS_38 => SharedReg145_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_39_cast,
                 iS_39 => SharedReg212_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_40_cast,
                 iS_4 => SharedReg28_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_5_cast,
                 iS_40 => SharedReg100_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_41_cast,
                 iS_41 => SharedReg274_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_42_cast,
                 iS_42 => SharedReg260_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_43_cast,
                 iS_43 => SharedReg153_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_44_cast,
                 iS_44 => SharedReg111_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_45_cast,
                 iS_45 => Delay871No_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_46_cast,
                 iS_46 => SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_47_cast,
                 iS_47 => SharedReg260_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_48_cast,
                 iS_48 => SharedReg87_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_49_cast,
                 iS_49 => SharedReg167_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_50_cast,
                 iS_5 => SharedReg107_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_6_cast,
                 iS_50 => SharedReg223_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_51_cast,
                 iS_51 => SharedReg274_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_52_cast,
                 iS_52 => SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_53_cast,
                 iS_53 => SharedReg162_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_54_cast,
                 iS_54 => SharedReg199_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_55_cast,
                 iS_55 => SharedReg264_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_56_cast,
                 iS_56 => SharedReg271_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_57_cast,
                 iS_57 => SharedReg272_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_58_cast,
                 iS_58 => SharedReg147_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_59_cast,
                 iS_6 => SharedReg256_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_7_cast,
                 iS_7 => SharedReg274_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_8_cast,
                 iS_8 => SharedReg274_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_9_cast,
                 iS_9 => SharedReg220_out_to_MUX_Sum10_3_impl_1_parent_implementedSystem_port_10_cast,
                 iSel => ModCount591_out,
                 oMux => MUX_Sum10_3_impl_1_out);

   Delay1No15_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => MUX_Sum10_3_impl_1_out,
                 Y => Delay1No15_out);
   Y_0_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Y_0_IEEE,
                 X => Delay1No16_out);
Y_0 <= Y_0_IEEE;

   Delay1No16_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg275_out,
                 Y => Delay1No16_out);
   Y_1_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Y_1_IEEE,
                 X => Delay1No17_out);
Y_1 <= Y_1_IEEE;

   Delay1No17_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg296_out,
                 Y => Delay1No17_out);
   Y_2_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Y_2_IEEE,
                 X => Delay1No18_out);
Y_2 <= Y_2_IEEE;

   Delay1No18_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg317_out,
                 Y => Delay1No18_out);
   Y_3_instance: OutputIEEE_8_23_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => Y_3_IEEE,
                 X => Delay1No19_out);
Y_3 <= Y_3_IEEE;

   Delay1No19_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg338_out,
                 Y => Delay1No19_out);

   Delay871No_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg55_out,
                 Y => Delay871No_out);

   Delay871No1_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg111_out,
                 Y => Delay871No1_out);

   Delay871No2_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg168_out,
                 Y => Delay871No2_out);

   Delay872No_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg225_out,
                 Y => Delay872No_out);

   Delay47No7_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg270_out,
                 Y => Delay47No7_out);

   Delay15No6_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg273_out,
                 Y => Delay15No6_out);

   Delay123No_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg295_out,
                 Y => Delay123No_out);

   Delay123No1_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg316_out,
                 Y => Delay123No1_out);

   Delay123No2_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg337_out,
                 Y => Delay123No2_out);

   Delay123No3_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg358_out,
                 Y => Delay123No3_out);

   MUX_Product_0_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product_0_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount591_out,
                 Output => MUX_Product_0_impl_0_LUT_out);

   MUX_Product_0_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product_0_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount591_out,
                 Output => MUX_Product_0_impl_1_LUT_out);

   MUX_Product_2_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product_2_impl_0_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount591_out,
                 Output => MUX_Product_2_impl_0_LUT_out);

   MUX_Product_2_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product_2_impl_1_LUT_wIn_6_wOut_6_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount591_out,
                 Output => MUX_Product_2_impl_1_LUT_out);

   MUX_Product1_2_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product1_2_impl_0_LUT_wIn_6_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount591_out,
                 Output => MUX_Product1_2_impl_0_LUT_out);

   MUX_Product1_2_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product1_2_impl_1_LUT_wIn_6_wOut_5_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount591_out,
                 Output => MUX_Product1_2_impl_1_LUT_out);

   MUX_Product10_3_impl_0_LUT_instance: GenericLut_LUTData_MUX_Product10_3_impl_0_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount591_out,
                 Output => MUX_Product10_3_impl_0_LUT_out);

   MUX_Product10_3_impl_1_LUT_instance: GenericLut_LUTData_MUX_Product10_3_impl_1_LUT_wIn_6_wOut_3_wrapper_component  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Input => ModCount591_out,
                 Output => MUX_Product10_3_impl_1_LUT_out);

   SharedReg_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => X_0_out,
                 Y => SharedReg_out);

   SharedReg1_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg_out,
                 Y => SharedReg1_out);

   SharedReg2_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg1_out,
                 Y => SharedReg2_out);

   SharedReg3_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg2_out,
                 Y => SharedReg3_out);

   SharedReg4_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg3_out,
                 Y => SharedReg4_out);

   SharedReg5_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg4_out,
                 Y => SharedReg5_out);

   SharedReg6_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg5_out,
                 Y => SharedReg6_out);

   SharedReg7_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg6_out,
                 Y => SharedReg7_out);

   SharedReg8_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg7_out,
                 Y => SharedReg8_out);

   SharedReg9_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg8_out,
                 Y => SharedReg9_out);

   SharedReg10_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg9_out,
                 Y => SharedReg10_out);

   SharedReg11_instance: Delay_34_DelayLength_28_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=28 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg10_out,
                 Y => SharedReg11_out);

   SharedReg12_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg11_out,
                 Y => SharedReg12_out);

   SharedReg13_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg12_out,
                 Y => SharedReg13_out);

   SharedReg14_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg13_out,
                 Y => SharedReg14_out);

   SharedReg15_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg14_out,
                 Y => SharedReg15_out);

   SharedReg16_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg15_out,
                 Y => SharedReg16_out);

   SharedReg17_instance: Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=38 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg16_out,
                 Y => SharedReg17_out);

   SharedReg18_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg17_out,
                 Y => SharedReg18_out);

   SharedReg19_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg18_out,
                 Y => SharedReg19_out);

   SharedReg20_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg19_out,
                 Y => SharedReg20_out);

   SharedReg21_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg20_out,
                 Y => SharedReg21_out);

   SharedReg22_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg21_out,
                 Y => SharedReg22_out);

   SharedReg23_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg22_out,
                 Y => SharedReg23_out);

   SharedReg24_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg23_out,
                 Y => SharedReg24_out);

   SharedReg25_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg24_out,
                 Y => SharedReg25_out);

   SharedReg26_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg25_out,
                 Y => SharedReg26_out);

   SharedReg27_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg26_out,
                 Y => SharedReg27_out);

   SharedReg28_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg27_out,
                 Y => SharedReg28_out);

   SharedReg29_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg28_out,
                 Y => SharedReg29_out);

   SharedReg30_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg29_out,
                 Y => SharedReg30_out);

   SharedReg31_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg30_out,
                 Y => SharedReg31_out);

   SharedReg32_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg31_out,
                 Y => SharedReg32_out);

   SharedReg33_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg32_out,
                 Y => SharedReg33_out);

   SharedReg34_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg33_out,
                 Y => SharedReg34_out);

   SharedReg35_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg34_out,
                 Y => SharedReg35_out);

   SharedReg36_instance: Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=38 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg35_out,
                 Y => SharedReg36_out);

   SharedReg37_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg36_out,
                 Y => SharedReg37_out);

   SharedReg38_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg37_out,
                 Y => SharedReg38_out);

   SharedReg39_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg38_out,
                 Y => SharedReg39_out);

   SharedReg40_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg39_out,
                 Y => SharedReg40_out);

   SharedReg41_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg40_out,
                 Y => SharedReg41_out);

   SharedReg42_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg41_out,
                 Y => SharedReg42_out);

   SharedReg43_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg42_out,
                 Y => SharedReg43_out);

   SharedReg44_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg43_out,
                 Y => SharedReg44_out);

   SharedReg45_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg44_out,
                 Y => SharedReg45_out);

   SharedReg46_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg45_out,
                 Y => SharedReg46_out);

   SharedReg47_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg46_out,
                 Y => SharedReg47_out);

   SharedReg48_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg47_out,
                 Y => SharedReg48_out);

   SharedReg49_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg48_out,
                 Y => SharedReg49_out);

   SharedReg50_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg49_out,
                 Y => SharedReg50_out);

   SharedReg51_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg50_out,
                 Y => SharedReg51_out);

   SharedReg52_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg51_out,
                 Y => SharedReg52_out);

   SharedReg53_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg52_out,
                 Y => SharedReg53_out);

   SharedReg54_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg53_out,
                 Y => SharedReg54_out);

   SharedReg55_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg54_out,
                 Y => SharedReg55_out);

   SharedReg56_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => X_1_out,
                 Y => SharedReg56_out);

   SharedReg57_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg56_out,
                 Y => SharedReg57_out);

   SharedReg58_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg57_out,
                 Y => SharedReg58_out);

   SharedReg59_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg58_out,
                 Y => SharedReg59_out);

   SharedReg60_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg59_out,
                 Y => SharedReg60_out);

   SharedReg61_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg60_out,
                 Y => SharedReg61_out);

   SharedReg62_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg61_out,
                 Y => SharedReg62_out);

   SharedReg63_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg62_out,
                 Y => SharedReg63_out);

   SharedReg64_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg63_out,
                 Y => SharedReg64_out);

   SharedReg65_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg64_out,
                 Y => SharedReg65_out);

   SharedReg66_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg65_out,
                 Y => SharedReg66_out);

   SharedReg67_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg66_out,
                 Y => SharedReg67_out);

   SharedReg68_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg67_out,
                 Y => SharedReg68_out);

   SharedReg69_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg68_out,
                 Y => SharedReg69_out);

   SharedReg70_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg69_out,
                 Y => SharedReg70_out);

   SharedReg71_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg70_out,
                 Y => SharedReg71_out);

   SharedReg72_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg71_out,
                 Y => SharedReg72_out);

   SharedReg73_instance: Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=38 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg72_out,
                 Y => SharedReg73_out);

   SharedReg74_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg73_out,
                 Y => SharedReg74_out);

   SharedReg75_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg74_out,
                 Y => SharedReg75_out);

   SharedReg76_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg75_out,
                 Y => SharedReg76_out);

   SharedReg77_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg76_out,
                 Y => SharedReg77_out);

   SharedReg78_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg77_out,
                 Y => SharedReg78_out);

   SharedReg79_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg78_out,
                 Y => SharedReg79_out);

   SharedReg80_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg79_out,
                 Y => SharedReg80_out);

   SharedReg81_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg80_out,
                 Y => SharedReg81_out);

   SharedReg82_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg81_out,
                 Y => SharedReg82_out);

   SharedReg83_instance: Delay_34_DelayLength_36_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=36 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg82_out,
                 Y => SharedReg83_out);

   SharedReg84_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg83_out,
                 Y => SharedReg84_out);

   SharedReg85_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg84_out,
                 Y => SharedReg85_out);

   SharedReg86_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg85_out,
                 Y => SharedReg86_out);

   SharedReg87_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg86_out,
                 Y => SharedReg87_out);

   SharedReg88_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg87_out,
                 Y => SharedReg88_out);

   SharedReg89_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg88_out,
                 Y => SharedReg89_out);

   SharedReg90_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg89_out,
                 Y => SharedReg90_out);

   SharedReg91_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg90_out,
                 Y => SharedReg91_out);

   SharedReg92_instance: Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=37 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg91_out,
                 Y => SharedReg92_out);

   SharedReg93_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg92_out,
                 Y => SharedReg93_out);

   SharedReg94_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg93_out,
                 Y => SharedReg94_out);

   SharedReg95_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg94_out,
                 Y => SharedReg95_out);

   SharedReg96_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg95_out,
                 Y => SharedReg96_out);

   SharedReg97_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg96_out,
                 Y => SharedReg97_out);

   SharedReg98_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg97_out,
                 Y => SharedReg98_out);

   SharedReg99_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg98_out,
                 Y => SharedReg99_out);

   SharedReg100_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg99_out,
                 Y => SharedReg100_out);

   SharedReg101_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg100_out,
                 Y => SharedReg101_out);

   SharedReg102_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg101_out,
                 Y => SharedReg102_out);

   SharedReg103_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg102_out,
                 Y => SharedReg103_out);

   SharedReg104_instance: Delay_34_DelayLength_8_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg103_out,
                 Y => SharedReg104_out);

   SharedReg105_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg104_out,
                 Y => SharedReg105_out);

   SharedReg106_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg105_out,
                 Y => SharedReg106_out);

   SharedReg107_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg106_out,
                 Y => SharedReg107_out);

   SharedReg108_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg107_out,
                 Y => SharedReg108_out);

   SharedReg109_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg108_out,
                 Y => SharedReg109_out);

   SharedReg110_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg109_out,
                 Y => SharedReg110_out);

   SharedReg111_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg110_out,
                 Y => SharedReg111_out);

   SharedReg112_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => X_2_out,
                 Y => SharedReg112_out);

   SharedReg113_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg112_out,
                 Y => SharedReg113_out);

   SharedReg114_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg113_out,
                 Y => SharedReg114_out);

   SharedReg115_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg114_out,
                 Y => SharedReg115_out);

   SharedReg116_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg115_out,
                 Y => SharedReg116_out);

   SharedReg117_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg116_out,
                 Y => SharedReg117_out);

   SharedReg118_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg117_out,
                 Y => SharedReg118_out);

   SharedReg119_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg118_out,
                 Y => SharedReg119_out);

   SharedReg120_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg119_out,
                 Y => SharedReg120_out);

   SharedReg121_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg120_out,
                 Y => SharedReg121_out);

   SharedReg122_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg121_out,
                 Y => SharedReg122_out);

   SharedReg123_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg122_out,
                 Y => SharedReg123_out);

   SharedReg124_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg123_out,
                 Y => SharedReg124_out);

   SharedReg125_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg124_out,
                 Y => SharedReg125_out);

   SharedReg126_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg125_out,
                 Y => SharedReg126_out);

   SharedReg127_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg126_out,
                 Y => SharedReg127_out);

   SharedReg128_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg127_out,
                 Y => SharedReg128_out);

   SharedReg129_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg128_out,
                 Y => SharedReg129_out);

   SharedReg130_instance: Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=38 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg129_out,
                 Y => SharedReg130_out);

   SharedReg131_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg130_out,
                 Y => SharedReg131_out);

   SharedReg132_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg131_out,
                 Y => SharedReg132_out);

   SharedReg133_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg132_out,
                 Y => SharedReg133_out);

   SharedReg134_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg133_out,
                 Y => SharedReg134_out);

   SharedReg135_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg134_out,
                 Y => SharedReg135_out);

   SharedReg136_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg135_out,
                 Y => SharedReg136_out);

   SharedReg137_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg136_out,
                 Y => SharedReg137_out);

   SharedReg138_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg137_out,
                 Y => SharedReg138_out);

   SharedReg139_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg138_out,
                 Y => SharedReg139_out);

   SharedReg140_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg139_out,
                 Y => SharedReg140_out);

   SharedReg141_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg140_out,
                 Y => SharedReg141_out);

   SharedReg142_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg141_out,
                 Y => SharedReg142_out);

   SharedReg143_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg142_out,
                 Y => SharedReg143_out);

   SharedReg144_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg143_out,
                 Y => SharedReg144_out);

   SharedReg145_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg144_out,
                 Y => SharedReg145_out);

   SharedReg146_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg145_out,
                 Y => SharedReg146_out);

   SharedReg147_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg146_out,
                 Y => SharedReg147_out);

   SharedReg148_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg147_out,
                 Y => SharedReg148_out);

   SharedReg149_instance: Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=37 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg148_out,
                 Y => SharedReg149_out);

   SharedReg150_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg149_out,
                 Y => SharedReg150_out);

   SharedReg151_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg150_out,
                 Y => SharedReg151_out);

   SharedReg152_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg151_out,
                 Y => SharedReg152_out);

   SharedReg153_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg152_out,
                 Y => SharedReg153_out);

   SharedReg154_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg153_out,
                 Y => SharedReg154_out);

   SharedReg155_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg154_out,
                 Y => SharedReg155_out);

   SharedReg156_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg155_out,
                 Y => SharedReg156_out);

   SharedReg157_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg156_out,
                 Y => SharedReg157_out);

   SharedReg158_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg157_out,
                 Y => SharedReg158_out);

   SharedReg159_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg158_out,
                 Y => SharedReg159_out);

   SharedReg160_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg159_out,
                 Y => SharedReg160_out);

   SharedReg161_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg160_out,
                 Y => SharedReg161_out);

   SharedReg162_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg161_out,
                 Y => SharedReg162_out);

   SharedReg163_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg162_out,
                 Y => SharedReg163_out);

   SharedReg164_instance: Delay_34_DelayLength_25_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=25 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg163_out,
                 Y => SharedReg164_out);

   SharedReg165_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg164_out,
                 Y => SharedReg165_out);

   SharedReg166_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg165_out,
                 Y => SharedReg166_out);

   SharedReg167_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg166_out,
                 Y => SharedReg167_out);

   SharedReg168_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg167_out,
                 Y => SharedReg168_out);

   SharedReg169_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => X_3_out,
                 Y => SharedReg169_out);

   SharedReg170_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg169_out,
                 Y => SharedReg170_out);

   SharedReg171_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg170_out,
                 Y => SharedReg171_out);

   SharedReg172_instance: Delay_34_DelayLength_16_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=16 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg171_out,
                 Y => SharedReg172_out);

   SharedReg173_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg172_out,
                 Y => SharedReg173_out);

   SharedReg174_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg173_out,
                 Y => SharedReg174_out);

   SharedReg175_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg174_out,
                 Y => SharedReg175_out);

   SharedReg176_instance: Delay_34_DelayLength_30_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=30 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg175_out,
                 Y => SharedReg176_out);

   SharedReg177_instance: Delay_34_DelayLength_24_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=24 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg176_out,
                 Y => SharedReg177_out);

   SharedReg178_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg177_out,
                 Y => SharedReg178_out);

   SharedReg179_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg178_out,
                 Y => SharedReg179_out);

   SharedReg180_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg179_out,
                 Y => SharedReg180_out);

   SharedReg181_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg180_out,
                 Y => SharedReg181_out);

   SharedReg182_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg181_out,
                 Y => SharedReg182_out);

   SharedReg183_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg182_out,
                 Y => SharedReg183_out);

   SharedReg184_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg183_out,
                 Y => SharedReg184_out);

   SharedReg185_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg184_out,
                 Y => SharedReg185_out);

   SharedReg186_instance: Delay_34_DelayLength_39_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=39 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg185_out,
                 Y => SharedReg186_out);

   SharedReg187_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg186_out,
                 Y => SharedReg187_out);

   SharedReg188_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg187_out,
                 Y => SharedReg188_out);

   SharedReg189_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg188_out,
                 Y => SharedReg189_out);

   SharedReg190_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg189_out,
                 Y => SharedReg190_out);

   SharedReg191_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg190_out,
                 Y => SharedReg191_out);

   SharedReg192_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg191_out,
                 Y => SharedReg192_out);

   SharedReg193_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg192_out,
                 Y => SharedReg193_out);

   SharedReg194_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg193_out,
                 Y => SharedReg194_out);

   SharedReg195_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg194_out,
                 Y => SharedReg195_out);

   SharedReg196_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg195_out,
                 Y => SharedReg196_out);

   SharedReg197_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg196_out,
                 Y => SharedReg197_out);

   SharedReg198_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg197_out,
                 Y => SharedReg198_out);

   SharedReg199_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg198_out,
                 Y => SharedReg199_out);

   SharedReg200_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg199_out,
                 Y => SharedReg200_out);

   SharedReg201_instance: Delay_34_DelayLength_19_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=19 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg200_out,
                 Y => SharedReg201_out);

   SharedReg202_instance: Delay_34_DelayLength_34_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=34 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg201_out,
                 Y => SharedReg202_out);

   SharedReg203_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg202_out,
                 Y => SharedReg203_out);

   SharedReg204_instance: Delay_34_DelayLength_18_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=18 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg203_out,
                 Y => SharedReg204_out);

   SharedReg205_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg204_out,
                 Y => SharedReg205_out);

   SharedReg206_instance: Delay_34_DelayLength_38_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=38 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg205_out,
                 Y => SharedReg206_out);

   SharedReg207_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg206_out,
                 Y => SharedReg207_out);

   SharedReg208_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg207_out,
                 Y => SharedReg208_out);

   SharedReg209_instance: Delay_34_DelayLength_21_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg208_out,
                 Y => SharedReg209_out);

   SharedReg210_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg209_out,
                 Y => SharedReg210_out);

   SharedReg211_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg210_out,
                 Y => SharedReg211_out);

   SharedReg212_instance: Delay_34_DelayLength_23_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=23 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg211_out,
                 Y => SharedReg212_out);

   SharedReg213_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg212_out,
                 Y => SharedReg213_out);

   SharedReg214_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg213_out,
                 Y => SharedReg214_out);

   SharedReg215_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg214_out,
                 Y => SharedReg215_out);

   SharedReg216_instance: Delay_34_DelayLength_13_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=13 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg215_out,
                 Y => SharedReg216_out);

   SharedReg217_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg216_out,
                 Y => SharedReg217_out);

   SharedReg218_instance: Delay_34_DelayLength_9_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=9 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg217_out,
                 Y => SharedReg218_out);

   SharedReg219_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg218_out,
                 Y => SharedReg219_out);

   SharedReg220_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg219_out,
                 Y => SharedReg220_out);

   SharedReg221_instance: Delay_34_DelayLength_26_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=26 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg220_out,
                 Y => SharedReg221_out);

   SharedReg222_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg221_out,
                 Y => SharedReg222_out);

   SharedReg223_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg222_out,
                 Y => SharedReg223_out);

   SharedReg224_instance: Delay_34_DelayLength_14_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=14 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg223_out,
                 Y => SharedReg224_out);

   SharedReg225_instance: Delay_34_DelayLength_10_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=10 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg224_out,
                 Y => SharedReg225_out);

   SharedReg226_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant_0_impl_out,
                 Y => SharedReg226_out);

   SharedReg227_instance: Delay_34_DelayLength_7_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=7 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant1_0_impl_out,
                 Y => SharedReg227_out);

   SharedReg228_instance: Delay_34_DelayLength_52_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=52 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant10_0_impl_out,
                 Y => SharedReg228_out);

   SharedReg229_instance: Delay_34_DelayLength_57_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=57 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant11_0_impl_out,
                 Y => SharedReg229_out);

   SharedReg230_instance: Delay_34_DelayLength_62_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=62 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant12_0_impl_out,
                 Y => SharedReg230_out);

   SharedReg231_instance: Delay_34_DelayLength_67_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=67 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant13_0_impl_out,
                 Y => SharedReg231_out);

   SharedReg232_instance: Delay_34_DelayLength_41_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=41 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant14_0_impl_out,
                 Y => SharedReg232_out);

   SharedReg233_instance: Delay_34_DelayLength_78_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=78 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant15_0_impl_out,
                 Y => SharedReg233_out);

   SharedReg234_instance: Delay_34_DelayLength_97_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=97 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant16_0_impl_out,
                 Y => SharedReg234_out);

   SharedReg235_instance: Delay_34_DelayLength_102_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=102 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant17_0_impl_out,
                 Y => SharedReg235_out);

   SharedReg236_instance: Delay_34_DelayLength_64_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=64 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant18_0_impl_out,
                 Y => SharedReg236_out);

   SharedReg237_instance: Delay_34_DelayLength_77_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=77 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant19_0_impl_out,
                 Y => SharedReg237_out);

   SharedReg238_instance: Delay_34_DelayLength_11_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=11 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant2_0_impl_out,
                 Y => SharedReg238_out);

   SharedReg239_instance: Delay_34_DelayLength_65_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=65 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant20_0_impl_out,
                 Y => SharedReg239_out);

   SharedReg240_instance: Delay_34_DelayLength_122_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=122 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant21_0_impl_out,
                 Y => SharedReg240_out);

   SharedReg241_instance: Delay_34_DelayLength_124_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=124 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant22_0_impl_out,
                 Y => SharedReg241_out);

   SharedReg242_instance: Delay_34_DelayLength_132_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=132 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant23_0_impl_out,
                 Y => SharedReg242_out);

   SharedReg243_instance: Delay_34_DelayLength_137_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=137 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant24_0_impl_out,
                 Y => SharedReg243_out);

   SharedReg244_instance: Delay_34_DelayLength_142_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=142 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant25_0_impl_out,
                 Y => SharedReg244_out);

   SharedReg245_instance: Delay_34_DelayLength_147_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=147 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant29_0_impl_out,
                 Y => SharedReg245_out);

   SharedReg246_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant3_0_impl_out,
                 Y => SharedReg246_out);

   SharedReg247_instance: Delay_34_DelayLength_107_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=107 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant32_0_impl_out,
                 Y => SharedReg247_out);

   SharedReg248_instance: Delay_34_DelayLength_99_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=99 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant33_0_impl_out,
                 Y => SharedReg248_out);

   SharedReg249_instance: Delay_34_DelayLength_104_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=104 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant34_0_impl_out,
                 Y => SharedReg249_out);

   SharedReg250_instance: Delay_34_DelayLength_20_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=20 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant4_0_impl_out,
                 Y => SharedReg250_out);

   SharedReg251_instance: Delay_34_DelayLength_27_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=27 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant5_0_impl_out,
                 Y => SharedReg251_out);

   SharedReg252_instance: Delay_34_DelayLength_32_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=32 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant6_0_impl_out,
                 Y => SharedReg252_out);

   SharedReg253_instance: Delay_34_DelayLength_37_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=37 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant7_0_impl_out,
                 Y => SharedReg253_out);

   SharedReg254_instance: Delay_34_DelayLength_42_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=42 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant8_0_impl_out,
                 Y => SharedReg254_out);

   SharedReg255_instance: Delay_34_DelayLength_47_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=47 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Constant9_0_impl_out,
                 Y => SharedReg255_out);

   SharedReg256_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product_0_impl_out,
                 Y => SharedReg256_out);

   SharedReg257_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg256_out,
                 Y => SharedReg257_out);

   SharedReg258_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg257_out,
                 Y => SharedReg258_out);

   SharedReg259_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg258_out,
                 Y => SharedReg259_out);

   SharedReg260_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg259_out,
                 Y => SharedReg260_out);

   SharedReg261_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg260_out,
                 Y => SharedReg261_out);

   SharedReg262_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg261_out,
                 Y => SharedReg262_out);

   SharedReg263_instance: Delay_34_DelayLength_29_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=29 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg262_out,
                 Y => SharedReg263_out);

   SharedReg264_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product_2_impl_out,
                 Y => SharedReg264_out);

   SharedReg265_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg264_out,
                 Y => SharedReg265_out);

   SharedReg266_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg265_out,
                 Y => SharedReg266_out);

   SharedReg267_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg266_out,
                 Y => SharedReg267_out);

   SharedReg268_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg267_out,
                 Y => SharedReg268_out);

   SharedReg269_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg268_out,
                 Y => SharedReg269_out);

   SharedReg270_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg269_out,
                 Y => SharedReg270_out);

   SharedReg271_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product1_2_impl_out,
                 Y => SharedReg271_out);

   SharedReg272_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg271_out,
                 Y => SharedReg272_out);

   SharedReg273_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg272_out,
                 Y => SharedReg273_out);

   SharedReg274_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Product10_3_impl_out,
                 Y => SharedReg274_out);

   SharedReg275_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Sum10_0_impl_out,
                 Y => SharedReg275_out);

   SharedReg276_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg275_out,
                 Y => SharedReg276_out);

   SharedReg277_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg276_out,
                 Y => SharedReg277_out);

   SharedReg278_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg277_out,
                 Y => SharedReg278_out);

   SharedReg279_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg278_out,
                 Y => SharedReg279_out);

   SharedReg280_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg279_out,
                 Y => SharedReg280_out);

   SharedReg281_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg280_out,
                 Y => SharedReg281_out);

   SharedReg282_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg281_out,
                 Y => SharedReg282_out);

   SharedReg283_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg282_out,
                 Y => SharedReg283_out);

   SharedReg284_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg283_out,
                 Y => SharedReg284_out);

   SharedReg285_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg284_out,
                 Y => SharedReg285_out);

   SharedReg286_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg285_out,
                 Y => SharedReg286_out);

   SharedReg287_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg286_out,
                 Y => SharedReg287_out);

   SharedReg288_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg287_out,
                 Y => SharedReg288_out);

   SharedReg289_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg288_out,
                 Y => SharedReg289_out);

   SharedReg290_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg289_out,
                 Y => SharedReg290_out);

   SharedReg291_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg290_out,
                 Y => SharedReg291_out);

   SharedReg292_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg291_out,
                 Y => SharedReg292_out);

   SharedReg293_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg292_out,
                 Y => SharedReg293_out);

   SharedReg294_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg293_out,
                 Y => SharedReg294_out);

   SharedReg295_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg294_out,
                 Y => SharedReg295_out);

   SharedReg296_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Sum10_1_impl_out,
                 Y => SharedReg296_out);

   SharedReg297_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg296_out,
                 Y => SharedReg297_out);

   SharedReg298_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg297_out,
                 Y => SharedReg298_out);

   SharedReg299_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg298_out,
                 Y => SharedReg299_out);

   SharedReg300_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg299_out,
                 Y => SharedReg300_out);

   SharedReg301_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg300_out,
                 Y => SharedReg301_out);

   SharedReg302_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg301_out,
                 Y => SharedReg302_out);

   SharedReg303_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg302_out,
                 Y => SharedReg303_out);

   SharedReg304_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg303_out,
                 Y => SharedReg304_out);

   SharedReg305_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg304_out,
                 Y => SharedReg305_out);

   SharedReg306_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg305_out,
                 Y => SharedReg306_out);

   SharedReg307_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg306_out,
                 Y => SharedReg307_out);

   SharedReg308_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg307_out,
                 Y => SharedReg308_out);

   SharedReg309_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg308_out,
                 Y => SharedReg309_out);

   SharedReg310_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg309_out,
                 Y => SharedReg310_out);

   SharedReg311_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg310_out,
                 Y => SharedReg311_out);

   SharedReg312_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg311_out,
                 Y => SharedReg312_out);

   SharedReg313_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg312_out,
                 Y => SharedReg313_out);

   SharedReg314_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg313_out,
                 Y => SharedReg314_out);

   SharedReg315_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg314_out,
                 Y => SharedReg315_out);

   SharedReg316_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg315_out,
                 Y => SharedReg316_out);

   SharedReg317_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Sum10_2_impl_out,
                 Y => SharedReg317_out);

   SharedReg318_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg317_out,
                 Y => SharedReg318_out);

   SharedReg319_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg318_out,
                 Y => SharedReg319_out);

   SharedReg320_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg319_out,
                 Y => SharedReg320_out);

   SharedReg321_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg320_out,
                 Y => SharedReg321_out);

   SharedReg322_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg321_out,
                 Y => SharedReg322_out);

   SharedReg323_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg322_out,
                 Y => SharedReg323_out);

   SharedReg324_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg323_out,
                 Y => SharedReg324_out);

   SharedReg325_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg324_out,
                 Y => SharedReg325_out);

   SharedReg326_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg325_out,
                 Y => SharedReg326_out);

   SharedReg327_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg326_out,
                 Y => SharedReg327_out);

   SharedReg328_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg327_out,
                 Y => SharedReg328_out);

   SharedReg329_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg328_out,
                 Y => SharedReg329_out);

   SharedReg330_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg329_out,
                 Y => SharedReg330_out);

   SharedReg331_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg330_out,
                 Y => SharedReg331_out);

   SharedReg332_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg331_out,
                 Y => SharedReg332_out);

   SharedReg333_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg332_out,
                 Y => SharedReg333_out);

   SharedReg334_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg333_out,
                 Y => SharedReg334_out);

   SharedReg335_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg334_out,
                 Y => SharedReg335_out);

   SharedReg336_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg335_out,
                 Y => SharedReg336_out);

   SharedReg337_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg336_out,
                 Y => SharedReg337_out);

   SharedReg338_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => Sum10_3_impl_out,
                 Y => SharedReg338_out);

   SharedReg339_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg338_out,
                 Y => SharedReg339_out);

   SharedReg340_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg339_out,
                 Y => SharedReg340_out);

   SharedReg341_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg340_out,
                 Y => SharedReg341_out);

   SharedReg342_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg341_out,
                 Y => SharedReg342_out);

   SharedReg343_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg342_out,
                 Y => SharedReg343_out);

   SharedReg344_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg343_out,
                 Y => SharedReg344_out);

   SharedReg345_instance: Delay_34_DelayLength_4_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=4 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg344_out,
                 Y => SharedReg345_out);

   SharedReg346_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg345_out,
                 Y => SharedReg346_out);

   SharedReg347_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg346_out,
                 Y => SharedReg347_out);

   SharedReg348_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg347_out,
                 Y => SharedReg348_out);

   SharedReg349_instance: Delay_34_DelayLength_2_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg348_out,
                 Y => SharedReg349_out);

   SharedReg350_instance: Delay_34_DelayLength_35_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=35 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg349_out,
                 Y => SharedReg350_out);

   SharedReg351_instance: Delay_34_DelayLength_1_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg350_out,
                 Y => SharedReg351_out);

   SharedReg352_instance: Delay_34_DelayLength_5_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg351_out,
                 Y => SharedReg352_out);

   SharedReg353_instance: Delay_34_DelayLength_15_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=15 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg352_out,
                 Y => SharedReg353_out);

   SharedReg354_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg353_out,
                 Y => SharedReg354_out);

   SharedReg355_instance: Delay_34_DelayLength_12_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=12 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg354_out,
                 Y => SharedReg355_out);

   SharedReg356_instance: Delay_34_DelayLength_6_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=6 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg355_out,
                 Y => SharedReg356_out);

   SharedReg357_instance: Delay_34_DelayLength_17_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=17 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg356_out,
                 Y => SharedReg357_out);

   SharedReg358_instance: Delay_34_DelayLength_3_initialCondition_0000000000000000000000000000000000_component  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => SharedReg357_out,
                 Y => SharedReg358_out);
end architecture;

